magic
tech scmos
timestamp 1554483974
<< m3contact >>
rect -2 -2 2 2
<< metal3 >>
rect -3 2 3 3
rect -3 -2 -2 2
rect 2 -2 3 2
rect -3 -3 3 -2
<< end >>
