magic
tech scmos
timestamp 1554483974
<< m2contact >>
rect -2 -2 2 2
<< end >>
