magic
tech scmos
timestamp 1522810115
<< nwell >>
rect 20 740 280 1000
rect 17 429 283 653
rect -3 249 303 330
rect -3 11 11 249
rect 289 11 303 249
rect -3 -3 303 11
<< pwell >>
rect -3 656 303 673
rect -3 426 14 656
rect 286 426 303 656
rect -3 340 303 426
rect 11 11 289 249
<< ptransistor >>
rect 38 626 138 629
rect 162 626 262 629
rect 38 582 138 585
rect 38 562 138 565
rect 162 582 262 585
rect 162 562 262 565
rect 38 518 138 521
rect 38 497 138 500
rect 162 518 262 521
rect 162 497 262 500
rect 38 453 138 456
rect 162 453 262 456
<< pdiffusion >>
rect 38 636 138 638
rect 38 632 41 636
rect 120 632 138 636
rect 38 629 138 632
rect 38 610 138 626
rect 38 601 56 610
rect 120 601 138 610
rect 38 585 138 601
rect 162 636 262 638
rect 162 632 180 636
rect 259 632 262 636
rect 162 629 262 632
rect 38 578 138 582
rect 38 569 41 578
rect 120 569 138 578
rect 38 565 138 569
rect 38 546 138 562
rect 38 537 56 546
rect 120 537 138 546
rect 38 521 138 537
rect 162 610 262 626
rect 162 601 180 610
rect 244 601 262 610
rect 162 585 262 601
rect 162 578 262 582
rect 162 569 180 578
rect 259 569 262 578
rect 162 565 262 569
rect 38 514 138 518
rect 38 510 41 514
rect 120 510 138 514
rect 38 508 138 510
rect 38 504 41 508
rect 120 504 138 508
rect 38 500 138 504
rect 38 481 138 497
rect 38 472 56 481
rect 120 472 138 481
rect 38 456 138 472
rect 162 546 262 562
rect 162 537 180 546
rect 244 537 262 546
rect 162 521 262 537
rect 162 514 262 518
rect 162 510 180 514
rect 259 510 262 514
rect 162 508 262 510
rect 162 504 180 508
rect 259 504 262 508
rect 162 500 262 504
rect 38 449 138 453
rect 38 445 41 449
rect 120 445 138 449
rect 38 444 138 445
rect 162 481 262 497
rect 162 472 180 481
rect 244 472 262 481
rect 162 456 262 472
rect 162 449 262 453
rect 162 445 180 449
rect 259 445 262 449
rect 162 444 262 445
<< pdcontact >>
rect 41 632 120 636
rect 56 601 120 610
rect 180 632 259 636
rect 41 569 120 578
rect 56 537 120 546
rect 180 601 244 610
rect 180 569 259 578
rect 41 510 120 514
rect 41 504 120 508
rect 56 472 120 481
rect 180 537 244 546
rect 180 510 259 514
rect 180 504 259 508
rect 41 445 120 449
rect 180 472 244 481
rect 180 445 259 449
<< psubstratepdiff >>
rect 0 669 300 670
rect 0 660 1 669
rect 130 660 170 669
rect 299 660 300 669
rect 0 659 300 660
rect 0 658 11 659
rect 0 424 1 658
rect 10 424 11 658
rect 289 658 300 659
rect 0 423 11 424
rect 289 424 290 658
rect 299 424 300 658
rect 289 423 300 424
rect 0 418 300 423
rect 0 414 3 418
rect 297 414 300 418
rect 0 408 300 414
rect 0 404 3 408
rect 297 404 300 408
rect 0 398 300 404
rect 0 394 3 398
rect 297 394 300 398
rect 0 388 300 394
rect 0 384 3 388
rect 297 384 300 388
rect 0 378 300 384
rect 0 374 3 378
rect 297 374 300 378
rect 0 368 300 374
rect 0 364 3 368
rect 297 364 300 368
rect 0 358 300 364
rect 0 354 3 358
rect 297 354 300 358
rect 0 348 300 354
rect 0 344 3 348
rect 297 344 300 348
rect 0 343 300 344
rect 14 245 286 246
rect 14 231 15 245
rect 284 231 286 245
rect 14 229 286 231
rect 14 225 15 229
rect 284 225 286 229
rect 14 219 286 225
rect 14 215 15 219
rect 284 215 286 219
rect 14 209 286 215
rect 14 205 15 209
rect 284 205 286 209
rect 14 199 286 205
rect 14 195 15 199
rect 284 195 286 199
rect 14 189 286 195
rect 14 185 15 189
rect 284 185 286 189
rect 14 179 286 185
rect 14 175 15 179
rect 284 175 286 179
rect 14 169 286 175
rect 14 165 15 169
rect 284 165 286 169
rect 14 159 286 165
rect 14 155 15 159
rect 284 155 286 159
rect 14 149 286 155
rect 14 145 15 149
rect 284 145 286 149
rect 14 139 286 145
rect 14 135 15 139
rect 284 135 286 139
rect 14 129 286 135
rect 14 125 15 129
rect 284 125 286 129
rect 14 119 286 125
rect 14 115 15 119
rect 284 115 286 119
rect 14 109 286 115
rect 14 105 15 109
rect 284 105 286 109
rect 14 99 286 105
rect 14 95 15 99
rect 284 95 286 99
rect 14 89 286 95
rect 14 85 15 89
rect 284 85 286 89
rect 14 79 286 85
rect 14 75 15 79
rect 284 75 286 79
rect 14 69 286 75
rect 14 65 15 69
rect 284 65 286 69
rect 14 59 286 65
rect 14 55 15 59
rect 284 55 286 59
rect 14 49 286 55
rect 14 45 15 49
rect 284 45 286 49
rect 14 39 286 45
rect 14 35 15 39
rect 284 35 286 39
rect 14 29 286 35
rect 14 25 15 29
rect 284 25 286 29
rect 14 19 286 25
rect 14 15 15 19
rect 284 15 286 19
rect 14 14 286 15
<< nsubstratendiff >>
rect 20 649 280 650
rect 20 445 26 649
rect 30 647 270 649
rect 30 643 36 647
rect 120 643 180 647
rect 264 643 270 647
rect 30 640 270 643
rect 36 638 138 640
rect 142 615 158 640
rect 162 638 264 640
rect 142 611 143 615
rect 157 611 158 615
rect 142 605 158 611
rect 142 601 143 605
rect 157 601 158 605
rect 142 595 158 601
rect 142 591 143 595
rect 157 591 158 595
rect 142 551 158 591
rect 142 547 143 551
rect 157 547 158 551
rect 142 541 158 547
rect 142 537 143 541
rect 157 537 158 541
rect 142 531 158 537
rect 142 527 143 531
rect 157 527 158 531
rect 142 486 158 527
rect 142 482 143 486
rect 157 482 158 486
rect 142 476 158 482
rect 142 472 143 476
rect 157 472 158 476
rect 142 466 158 472
rect 142 462 143 466
rect 157 462 158 466
rect 20 442 30 445
rect 38 442 138 444
rect 142 442 158 462
rect 162 442 262 444
rect 274 445 280 649
rect 270 442 280 445
rect 20 441 280 442
rect 20 432 21 441
rect 120 432 180 441
rect 279 432 280 441
rect 0 326 300 327
rect 0 322 2 326
rect 96 322 143 326
rect 157 322 204 326
rect 298 322 300 326
rect 0 316 300 322
rect 0 312 2 316
rect 96 312 143 316
rect 157 312 204 316
rect 298 312 300 316
rect 0 306 300 312
rect 0 302 2 306
rect 96 302 143 306
rect 157 302 204 306
rect 298 302 300 306
rect 0 296 300 302
rect 0 292 2 296
rect 96 292 143 296
rect 157 292 204 296
rect 298 292 300 296
rect 0 286 300 292
rect 0 282 2 286
rect 96 282 143 286
rect 157 282 204 286
rect 298 282 300 286
rect 0 276 300 282
rect 0 272 2 276
rect 96 272 143 276
rect 157 272 204 276
rect 298 272 300 276
rect 0 266 300 272
rect 0 262 2 266
rect 96 262 143 266
rect 157 262 204 266
rect 298 262 300 266
rect 0 256 300 262
rect 0 2 2 256
rect 6 8 8 256
rect 97 252 143 256
rect 157 252 203 256
rect 292 8 294 256
rect 6 6 294 8
rect 6 2 10 6
rect 94 2 206 6
rect 290 2 294 6
rect 298 2 300 256
rect 0 0 300 2
<< psubstratepcontact >>
rect 1 660 130 669
rect 170 660 299 669
rect 1 424 10 658
rect 290 424 299 658
rect 3 414 297 418
rect 3 404 297 408
rect 3 394 297 398
rect 3 384 297 388
rect 3 374 297 378
rect 3 364 297 368
rect 3 354 297 358
rect 3 344 297 348
rect 15 231 284 245
rect 15 225 284 229
rect 15 215 284 219
rect 15 205 284 209
rect 15 195 284 199
rect 15 185 284 189
rect 15 175 284 179
rect 15 165 284 169
rect 15 155 284 159
rect 15 145 284 149
rect 15 135 284 139
rect 15 125 284 129
rect 15 115 284 119
rect 15 105 284 109
rect 15 95 284 99
rect 15 85 284 89
rect 15 75 284 79
rect 15 65 284 69
rect 15 55 284 59
rect 15 45 284 49
rect 15 35 284 39
rect 15 25 284 29
rect 15 15 284 19
<< nsubstratencontact >>
rect 26 445 30 649
rect 36 643 120 647
rect 180 643 264 647
rect 143 611 157 615
rect 143 601 157 605
rect 143 591 157 595
rect 143 547 157 551
rect 143 537 157 541
rect 143 527 157 531
rect 143 482 157 486
rect 143 472 157 476
rect 143 462 157 466
rect 270 445 274 649
rect 21 432 120 441
rect 180 432 279 441
rect 2 322 96 326
rect 143 322 157 326
rect 204 322 298 326
rect 2 312 96 316
rect 143 312 157 316
rect 204 312 298 316
rect 2 302 96 306
rect 143 302 157 306
rect 204 302 298 306
rect 2 292 96 296
rect 143 292 157 296
rect 204 292 298 296
rect 2 282 96 286
rect 143 282 157 286
rect 204 282 298 286
rect 2 272 96 276
rect 143 272 157 276
rect 204 272 298 276
rect 2 262 96 266
rect 143 262 157 266
rect 204 262 298 266
rect 2 2 6 256
rect 8 252 97 256
rect 143 252 157 256
rect 203 252 292 256
rect 10 2 94 6
rect 206 2 290 6
rect 294 2 298 256
<< polysilicon >>
rect 2 715 17 718
rect 20 715 35 718
rect 8 703 11 715
rect 20 712 23 715
rect 32 712 35 715
rect 20 709 35 712
rect 20 703 23 709
rect 32 703 35 709
rect 38 715 41 718
rect 38 712 47 715
rect 38 703 41 712
rect 44 709 47 712
rect 50 709 53 718
rect 44 706 53 709
rect 50 703 53 706
rect 56 715 59 718
rect 56 712 65 715
rect 56 703 59 712
rect 62 709 65 712
rect 68 709 71 718
rect 62 706 71 709
rect 68 703 71 706
rect 74 715 89 718
rect 92 715 107 718
rect 74 712 77 715
rect 92 712 95 715
rect 104 712 107 715
rect 74 709 89 712
rect 92 709 107 712
rect 74 706 77 709
rect 74 703 89 706
rect 92 703 95 709
rect 101 703 104 709
rect 194 707 209 710
rect 194 695 197 707
rect 200 701 203 707
rect 206 695 209 707
rect 212 707 227 710
rect 212 698 215 707
rect 224 698 227 707
rect 230 707 245 710
rect 248 707 263 710
rect 266 707 281 710
rect 230 704 233 707
rect 230 701 245 704
rect 242 698 245 701
rect 254 698 257 707
rect 266 704 269 707
rect 266 701 281 704
rect 278 698 281 701
rect 212 695 227 698
rect 230 695 245 698
rect 248 695 263 698
rect 266 695 281 698
rect 42 689 57 692
rect 60 689 75 692
rect 78 689 93 692
rect 42 680 45 689
rect 60 686 63 689
rect 78 686 81 689
rect 60 683 75 686
rect 78 683 93 686
rect 60 680 63 683
rect 90 680 93 683
rect 42 677 57 680
rect 60 677 75 680
rect 78 677 93 680
rect 31 626 38 629
rect 138 626 140 629
rect 31 457 32 626
rect 36 585 37 626
rect 160 626 162 629
rect 262 626 269 629
rect 36 582 38 585
rect 138 582 140 585
rect 36 565 37 582
rect 36 562 38 565
rect 138 562 140 565
rect 36 521 37 562
rect 263 585 264 626
rect 160 582 162 585
rect 262 582 264 585
rect 263 565 264 582
rect 160 562 162 565
rect 262 562 264 565
rect 36 518 38 521
rect 138 518 140 521
rect 36 500 37 518
rect 36 497 38 500
rect 138 497 140 500
rect 36 457 37 497
rect 31 456 37 457
rect 263 521 264 562
rect 160 518 162 521
rect 262 518 264 521
rect 263 500 264 518
rect 160 497 162 500
rect 262 497 264 500
rect 31 453 38 456
rect 138 453 140 456
rect 263 457 264 497
rect 268 457 269 626
rect 263 456 269 457
rect 160 453 162 456
rect 262 453 269 456
<< polycontact >>
rect 32 457 36 626
rect 264 457 268 626
<< metal1 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 62 730 238 740
rect 72 720 228 730
rect 82 710 218 720
rect 92 700 208 710
rect 102 670 198 700
rect 0 669 300 670
rect 0 660 1 669
rect 130 660 170 669
rect 299 660 300 669
rect 0 659 300 660
rect 0 658 11 659
rect 0 424 1 658
rect 10 424 11 658
rect 102 653 198 659
rect 289 658 300 659
rect 36 649 120 650
rect 20 445 21 649
rect 25 445 26 649
rect 30 647 120 649
rect 30 643 36 647
rect 30 642 120 643
rect 30 638 36 642
rect 30 636 120 638
rect 30 632 41 636
rect 30 626 120 632
rect 30 457 32 626
rect 36 625 120 626
rect 36 586 39 625
rect 48 621 52 625
rect 116 621 120 625
rect 48 590 51 621
rect 123 618 177 653
rect 180 649 280 650
rect 180 647 270 649
rect 264 643 270 647
rect 180 642 270 643
rect 264 638 270 642
rect 180 636 270 638
rect 259 632 270 636
rect 180 626 270 632
rect 180 625 264 626
rect 180 621 184 625
rect 248 621 252 625
rect 56 610 140 618
rect 120 601 140 610
rect 56 593 140 601
rect 48 586 52 590
rect 116 586 120 590
rect 36 578 120 586
rect 36 569 41 578
rect 36 561 120 569
rect 36 522 39 561
rect 48 557 52 561
rect 116 557 120 561
rect 123 588 140 593
rect 143 610 157 611
rect 143 605 157 606
rect 143 600 157 601
rect 143 595 157 596
rect 160 610 244 618
rect 160 601 180 610
rect 160 593 244 601
rect 160 588 177 593
rect 249 590 252 621
rect 48 526 51 557
rect 123 554 177 588
rect 180 586 184 590
rect 248 586 252 590
rect 261 586 264 625
rect 180 578 264 586
rect 259 569 264 578
rect 180 561 264 569
rect 180 557 184 561
rect 248 557 252 561
rect 56 546 140 554
rect 120 537 140 546
rect 56 529 140 537
rect 48 522 52 526
rect 116 522 120 526
rect 36 514 120 522
rect 36 510 41 514
rect 36 508 120 510
rect 36 504 41 508
rect 36 496 120 504
rect 36 457 39 496
rect 48 492 52 496
rect 116 492 120 496
rect 123 524 140 529
rect 143 546 157 547
rect 143 541 157 542
rect 143 536 157 537
rect 143 531 157 532
rect 160 546 244 554
rect 160 537 180 546
rect 160 529 244 537
rect 160 524 177 529
rect 249 526 252 557
rect 48 461 51 492
rect 123 489 177 524
rect 180 522 184 526
rect 248 522 252 526
rect 261 522 264 561
rect 180 514 264 522
rect 259 510 264 514
rect 180 508 264 510
rect 259 504 264 508
rect 180 496 264 504
rect 180 492 184 496
rect 248 492 252 496
rect 56 481 140 489
rect 120 472 140 481
rect 56 464 140 472
rect 48 457 52 461
rect 116 457 120 461
rect 30 449 120 457
rect 30 445 41 449
rect 20 441 120 445
rect 20 432 21 441
rect 123 459 140 464
rect 143 481 157 482
rect 143 476 157 477
rect 143 471 157 472
rect 143 466 157 467
rect 160 481 244 489
rect 160 472 180 481
rect 160 464 244 472
rect 160 459 177 464
rect 249 461 252 492
rect 123 429 177 459
rect 180 457 184 461
rect 248 457 252 461
rect 261 457 264 496
rect 268 457 270 626
rect 180 449 270 457
rect 259 445 270 449
rect 274 445 275 649
rect 279 445 280 649
rect 180 441 280 445
rect 279 432 280 441
rect 0 423 11 424
rect 102 423 198 429
rect 289 424 290 658
rect 299 424 300 658
rect 289 423 300 424
rect 0 418 300 423
rect 0 414 3 418
rect 297 414 300 418
rect 0 413 300 414
rect 0 409 3 413
rect 297 409 300 413
rect 0 408 300 409
rect 0 404 3 408
rect 297 404 300 408
rect 0 403 300 404
rect 0 399 3 403
rect 297 399 300 403
rect 0 398 300 399
rect 0 394 3 398
rect 297 394 300 398
rect 0 393 300 394
rect 0 389 3 393
rect 297 389 300 393
rect 0 388 300 389
rect 0 384 3 388
rect 297 384 300 388
rect 0 383 300 384
rect 0 379 3 383
rect 297 379 300 383
rect 0 378 300 379
rect 0 374 3 378
rect 297 374 300 378
rect 0 373 300 374
rect 0 369 3 373
rect 297 369 300 373
rect 0 368 300 369
rect 0 364 3 368
rect 297 364 300 368
rect 0 363 300 364
rect 0 359 3 363
rect 297 359 300 363
rect 0 358 300 359
rect 0 354 3 358
rect 297 354 300 358
rect 0 353 300 354
rect 0 349 3 353
rect 297 349 300 353
rect 0 348 300 349
rect 0 344 3 348
rect 297 344 300 348
rect 102 329 198 344
rect 0 322 2 326
rect 96 322 99 326
rect 0 321 99 322
rect 0 317 2 321
rect 96 317 99 321
rect 0 316 99 317
rect 0 312 2 316
rect 96 312 99 316
rect 0 311 99 312
rect 0 307 2 311
rect 96 307 99 311
rect 0 306 99 307
rect 0 302 2 306
rect 96 302 99 306
rect 0 301 99 302
rect 0 297 2 301
rect 96 297 99 301
rect 0 296 99 297
rect 0 292 2 296
rect 96 292 99 296
rect 0 291 99 292
rect 0 287 2 291
rect 96 287 99 291
rect 0 286 99 287
rect 0 282 2 286
rect 96 282 99 286
rect 0 281 99 282
rect 0 277 2 281
rect 96 277 99 281
rect 0 276 99 277
rect 0 272 2 276
rect 96 272 99 276
rect 0 271 99 272
rect 0 267 2 271
rect 96 267 99 271
rect 0 266 99 267
rect 0 262 2 266
rect 96 262 99 266
rect 0 261 99 262
rect 0 257 7 261
rect 96 257 99 261
rect 0 256 99 257
rect 0 2 2 256
rect 6 252 8 256
rect 97 252 99 256
rect 6 7 7 252
rect 102 246 140 329
rect 143 321 157 322
rect 143 316 157 317
rect 143 311 157 312
rect 143 306 157 307
rect 143 301 157 302
rect 143 296 157 297
rect 143 291 157 292
rect 143 286 157 287
rect 143 281 157 282
rect 143 276 157 277
rect 143 271 157 272
rect 143 266 157 267
rect 143 261 157 262
rect 143 256 157 257
rect 160 246 198 329
rect 201 322 204 326
rect 298 322 300 326
rect 201 321 300 322
rect 201 317 204 321
rect 298 317 300 321
rect 201 316 300 317
rect 201 312 204 316
rect 298 312 300 316
rect 201 311 300 312
rect 201 307 204 311
rect 298 307 300 311
rect 201 306 300 307
rect 201 302 204 306
rect 298 302 300 306
rect 201 301 300 302
rect 201 297 204 301
rect 298 297 300 301
rect 201 296 300 297
rect 201 292 204 296
rect 298 292 300 296
rect 201 291 300 292
rect 201 287 204 291
rect 298 287 300 291
rect 201 286 300 287
rect 201 282 204 286
rect 298 282 300 286
rect 201 281 300 282
rect 201 277 204 281
rect 298 277 300 281
rect 201 276 300 277
rect 201 272 204 276
rect 298 272 300 276
rect 201 271 300 272
rect 201 267 204 271
rect 298 267 300 271
rect 201 266 300 267
rect 201 262 204 266
rect 298 262 300 266
rect 201 261 300 262
rect 201 257 203 261
rect 292 257 300 261
rect 201 256 300 257
rect 201 252 203 256
rect 292 252 294 256
rect 102 245 198 246
rect 284 231 285 245
rect 15 229 285 231
rect 284 225 285 229
rect 15 224 285 225
rect 284 220 285 224
rect 15 219 285 220
rect 284 215 285 219
rect 15 214 285 215
rect 284 210 285 214
rect 15 209 285 210
rect 284 205 285 209
rect 15 204 285 205
rect 284 200 285 204
rect 15 199 285 200
rect 284 195 285 199
rect 15 194 285 195
rect 284 190 285 194
rect 15 189 285 190
rect 284 185 285 189
rect 15 184 285 185
rect 284 180 285 184
rect 15 179 285 180
rect 284 175 285 179
rect 15 174 285 175
rect 284 170 285 174
rect 15 169 285 170
rect 284 165 285 169
rect 15 164 285 165
rect 284 160 285 164
rect 15 159 285 160
rect 284 155 285 159
rect 15 154 285 155
rect 284 150 285 154
rect 15 149 285 150
rect 284 145 285 149
rect 15 144 285 145
rect 284 140 285 144
rect 15 139 285 140
rect 284 135 285 139
rect 15 134 285 135
rect 284 130 285 134
rect 15 129 285 130
rect 284 125 285 129
rect 15 124 285 125
rect 284 120 285 124
rect 15 119 285 120
rect 284 115 285 119
rect 15 114 285 115
rect 284 110 285 114
rect 15 109 285 110
rect 284 105 285 109
rect 15 104 285 105
rect 284 100 285 104
rect 15 99 285 100
rect 284 95 285 99
rect 15 94 285 95
rect 284 90 285 94
rect 15 89 285 90
rect 284 85 285 89
rect 15 84 285 85
rect 284 80 285 84
rect 15 79 285 80
rect 284 75 285 79
rect 15 74 285 75
rect 284 70 285 74
rect 15 69 285 70
rect 284 65 285 69
rect 15 64 285 65
rect 284 60 285 64
rect 15 59 285 60
rect 284 55 285 59
rect 15 54 285 55
rect 284 50 285 54
rect 15 49 285 50
rect 284 45 285 49
rect 15 44 285 45
rect 284 40 285 44
rect 15 39 285 40
rect 284 35 285 39
rect 15 34 285 35
rect 284 30 285 34
rect 15 29 285 30
rect 284 25 285 29
rect 15 24 285 25
rect 284 20 285 24
rect 15 19 285 20
rect 284 15 285 19
rect 6 6 99 7
rect 6 2 10 6
rect 94 2 99 6
rect 0 1 99 2
rect 102 6 198 15
rect 293 7 294 252
rect 102 2 103 6
rect 197 2 198 6
rect 102 -11 198 2
rect 201 6 294 7
rect 201 2 206 6
rect 290 2 294 6
rect 298 2 300 256
rect 201 1 300 2
<< m2contact >>
rect 21 445 25 649
rect 36 638 120 642
rect 39 586 48 625
rect 52 621 116 625
rect 180 638 264 642
rect 184 621 248 625
rect 52 586 116 590
rect 39 522 48 561
rect 52 557 116 561
rect 143 606 157 610
rect 143 596 157 600
rect 184 586 248 590
rect 252 586 261 625
rect 184 557 248 561
rect 52 522 116 526
rect 39 457 48 496
rect 52 492 116 496
rect 143 542 157 546
rect 143 532 157 536
rect 184 522 248 526
rect 252 522 261 561
rect 184 492 248 496
rect 52 457 116 461
rect 143 477 157 481
rect 143 467 157 471
rect 184 457 248 461
rect 252 457 261 496
rect 275 445 279 649
rect 3 409 297 413
rect 3 399 297 403
rect 3 389 297 393
rect 3 379 297 383
rect 3 369 297 373
rect 3 359 297 363
rect 3 349 297 353
rect 2 317 96 321
rect 2 307 96 311
rect 2 297 96 301
rect 2 287 96 291
rect 2 277 96 281
rect 2 267 96 271
rect 7 257 96 261
rect 143 317 157 321
rect 143 307 157 311
rect 143 297 157 301
rect 143 287 157 291
rect 143 277 157 281
rect 143 267 157 271
rect 143 257 157 261
rect 204 317 298 321
rect 204 307 298 311
rect 204 297 298 301
rect 204 287 298 291
rect 204 277 298 281
rect 204 267 298 271
rect 203 257 292 261
rect 15 220 284 224
rect 15 210 284 214
rect 15 200 284 204
rect 15 190 284 194
rect 15 180 284 184
rect 15 170 284 174
rect 15 160 284 164
rect 15 150 284 154
rect 15 140 284 144
rect 15 130 284 134
rect 15 120 284 124
rect 15 110 284 114
rect 15 100 284 104
rect 15 90 284 94
rect 15 80 284 84
rect 15 70 284 74
rect 15 60 284 64
rect 15 50 284 54
rect 15 40 284 44
rect 15 30 284 34
rect 15 20 284 24
rect 103 2 197 6
<< metal2 >>
rect 20 997 280 1000
rect 20 743 23 997
rect 277 743 280 997
rect 20 740 280 743
rect 0 649 300 670
rect 0 445 21 649
rect 25 642 275 649
rect 25 638 36 642
rect 120 638 180 642
rect 264 638 275 642
rect 25 625 275 638
rect 25 586 39 625
rect 48 621 52 625
rect 116 621 184 625
rect 248 621 252 625
rect 48 610 252 621
rect 48 606 143 610
rect 157 606 252 610
rect 48 600 252 606
rect 48 596 143 600
rect 157 596 252 600
rect 48 590 252 596
rect 48 586 52 590
rect 116 586 184 590
rect 248 586 252 590
rect 261 586 275 625
rect 25 561 275 586
rect 25 522 39 561
rect 48 557 52 561
rect 116 557 184 561
rect 248 557 252 561
rect 48 546 252 557
rect 48 542 143 546
rect 157 542 252 546
rect 48 536 252 542
rect 48 532 143 536
rect 157 532 252 536
rect 48 526 252 532
rect 48 522 52 526
rect 116 522 184 526
rect 248 522 252 526
rect 261 522 275 561
rect 25 496 275 522
rect 25 457 39 496
rect 48 492 52 496
rect 116 492 184 496
rect 248 492 252 496
rect 48 481 252 492
rect 48 477 143 481
rect 157 477 252 481
rect 48 471 252 477
rect 48 467 143 471
rect 157 467 252 471
rect 48 461 252 467
rect 48 457 52 461
rect 116 457 184 461
rect 248 457 252 461
rect 261 457 275 496
rect 25 445 275 457
rect 279 445 300 649
rect 0 440 300 445
rect 0 413 300 424
rect 0 409 3 413
rect 297 409 300 413
rect 0 403 300 409
rect 0 399 3 403
rect 297 399 300 403
rect 0 393 300 399
rect 0 389 3 393
rect 297 389 300 393
rect 0 383 300 389
rect 0 379 3 383
rect 297 379 300 383
rect 0 373 300 379
rect 0 369 3 373
rect 297 369 300 373
rect 0 363 300 369
rect 0 359 3 363
rect 297 359 300 363
rect 0 353 300 359
rect 0 349 3 353
rect 297 349 300 353
rect 0 344 300 349
rect 0 321 300 326
rect 0 317 2 321
rect 96 317 143 321
rect 157 317 204 321
rect 298 317 300 321
rect 0 311 300 317
rect 0 307 2 311
rect 96 307 143 311
rect 157 307 204 311
rect 298 307 300 311
rect 0 301 300 307
rect 0 297 2 301
rect 96 297 143 301
rect 157 297 204 301
rect 298 297 300 301
rect 0 291 300 297
rect 0 287 2 291
rect 96 287 143 291
rect 157 287 204 291
rect 298 287 300 291
rect 0 281 300 287
rect 0 277 2 281
rect 96 277 143 281
rect 157 277 204 281
rect 298 277 300 281
rect 0 271 300 277
rect 0 267 2 271
rect 96 267 143 271
rect 157 267 204 271
rect 298 267 300 271
rect 0 261 300 267
rect 0 257 7 261
rect 96 257 143 261
rect 157 257 203 261
rect 292 257 300 261
rect 0 246 300 257
rect 0 224 300 230
rect 0 220 15 224
rect 284 220 300 224
rect 0 214 300 220
rect 0 210 15 214
rect 284 210 300 214
rect 0 204 300 210
rect 0 200 15 204
rect 284 200 300 204
rect 0 194 300 200
rect 0 190 15 194
rect 284 190 300 194
rect 0 184 300 190
rect 0 180 15 184
rect 284 180 300 184
rect 0 174 300 180
rect 0 170 15 174
rect 284 170 300 174
rect 0 164 300 170
rect 0 160 15 164
rect 284 160 300 164
rect 0 154 300 160
rect 0 150 15 154
rect 284 150 300 154
rect 0 144 300 150
rect 0 140 15 144
rect 284 140 300 144
rect 0 134 300 140
rect 0 130 15 134
rect 284 130 300 134
rect 0 124 300 130
rect 0 120 15 124
rect 284 120 300 124
rect 0 114 300 120
rect 0 110 15 114
rect 284 110 300 114
rect 0 104 300 110
rect 0 100 15 104
rect 284 100 300 104
rect 0 94 300 100
rect 0 90 15 94
rect 284 90 300 94
rect 0 84 300 90
rect 0 80 15 84
rect 284 80 300 84
rect 0 74 300 80
rect 0 70 15 74
rect 284 70 300 74
rect 0 64 300 70
rect 0 60 15 64
rect 284 60 300 64
rect 0 54 300 60
rect 0 50 15 54
rect 284 50 300 54
rect 0 44 300 50
rect 0 40 15 44
rect 284 40 300 44
rect 0 34 300 40
rect 0 30 15 34
rect 284 30 300 34
rect 0 24 300 30
rect 0 20 15 24
rect 284 20 300 24
rect 0 6 300 20
rect 0 2 103 6
rect 197 2 300 6
rect 0 0 300 2
<< pad >>
rect 23 743 277 997
<< labels >>
rlabel metal1 150 0 150 0 8 GND!
rlabel metal2 132 540 132 540 6 vdd:2
rlabel metal1 150 -8 150 -8 1 GND!
<< end >>
