magic
tech scmos
timestamp 1553978028
<< nwell >>
rect -9 48 45 105
<< ntransistor >>
rect 7 6 9 26
rect 15 6 17 26
rect 23 6 25 26
rect 31 6 33 26
<< ptransistor >>
rect 7 54 9 94
rect 15 54 17 94
rect 23 54 25 94
rect 31 54 33 94
<< ndiffusion >>
rect 2 25 7 26
rect 6 6 7 25
rect 9 25 15 26
rect 9 6 10 25
rect 14 6 15 25
rect 17 25 23 26
rect 17 6 18 25
rect 22 6 23 25
rect 25 25 31 26
rect 25 6 26 25
rect 30 6 31 25
rect 33 25 38 26
rect 33 6 34 25
<< pdiffusion >>
rect 2 93 7 94
rect 6 54 7 93
rect 9 93 15 94
rect 9 54 10 93
rect 14 54 15 93
rect 17 93 23 94
rect 17 54 18 93
rect 22 54 23 93
rect 25 93 31 94
rect 25 54 26 93
rect 30 54 31 93
rect 33 93 38 94
rect 33 54 34 93
<< ndcontact >>
rect 2 6 6 25
rect 10 6 14 25
rect 18 6 22 25
rect 26 6 30 25
rect 34 6 38 25
<< pdcontact >>
rect 2 54 6 93
rect 10 54 14 93
rect 18 54 22 93
rect 26 54 30 93
rect 34 54 38 93
<< psubstratepcontact >>
rect -2 -2 2 2
rect 14 -2 18 2
rect 30 -2 34 2
<< nsubstratencontact >>
rect -2 98 2 102
rect 14 98 18 102
rect 30 98 34 102
<< polysilicon >>
rect 7 94 9 96
rect 15 94 17 96
rect 23 94 25 96
rect 31 94 33 96
rect 7 53 9 54
rect 15 53 17 54
rect 23 53 25 54
rect 31 53 33 54
rect 7 51 33 53
rect 7 33 9 51
rect 6 30 9 33
rect 6 29 33 30
rect 7 28 33 29
rect 7 26 9 28
rect 15 26 17 28
rect 23 26 25 28
rect 31 26 33 28
rect 7 4 9 6
rect 15 4 17 6
rect 23 4 25 6
rect 31 4 33 6
<< polycontact >>
rect 2 29 6 33
<< metal1 >>
rect -2 102 42 103
rect 2 98 14 102
rect 18 98 30 102
rect 34 98 42 102
rect -2 97 42 98
rect 2 93 6 97
rect 10 93 14 94
rect 18 93 22 97
rect 26 93 30 94
rect 34 93 38 97
rect 10 51 14 54
rect 26 51 30 54
rect 10 47 30 51
rect 2 33 6 37
rect 26 33 30 47
rect 10 29 30 33
rect 2 25 6 26
rect 10 25 14 29
rect 18 25 22 26
rect 26 25 30 29
rect 34 25 38 26
rect 2 3 6 6
rect 18 3 22 6
rect 34 3 38 6
rect -2 2 42 3
rect 2 -2 14 2
rect 18 -2 30 2
rect 34 -2 42 2
rect -2 -3 42 -2
<< m1p >>
rect 26 43 30 47
rect 2 33 6 37
<< labels >>
rlabel metal1 4 100 4 100 4 vdd
rlabel metal1 4 0 4 0 4 gnd
rlabel metal1 4 35 4 35 4 A
rlabel metal1 28 45 28 45 4 Y
<< end >>
