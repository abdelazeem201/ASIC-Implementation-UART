magic
tech scmos
timestamp 1555511723
<< polysilicon >>
rect 1 4033 291 4991
rect 336 4691 996 4997
rect 4010 4689 4694 4998
rect 4701 4965 4993 5000
rect 4701 4010 4991 4965
rect 1435 3354 2257 3661
rect 3477 2662 3621 3277
rect 1315 1207 1488 2043
rect 2823 1154 3318 1581
rect 2 256 308 992
rect 4700 263 4994 972
rect 4699 258 4994 263
rect 2 1 1005 256
rect 4009 3 4994 258
<< metal1 >>
rect 1029 3975 1139 3981
rect 1133 3923 1139 3975
rect 1323 3923 1329 3975
rect 1623 3923 1629 3975
rect 1923 3923 1929 3975
rect 2223 3923 2229 3975
rect 2523 3923 2529 3975
rect 1133 3917 2694 3923
rect 1133 2699 1139 3917
rect 1174 3744 1318 3750
rect 1312 3429 1318 3744
rect 2688 3493 2694 3917
rect 3123 3493 3129 3975
rect 3423 3503 3429 3975
rect 3723 3911 3729 3975
rect 3723 3905 3858 3911
rect 3852 3756 3858 3905
rect 3852 3729 3859 3756
rect 3852 3723 3975 3729
rect 3852 3666 3859 3723
rect 3423 3493 3428 3503
rect 2688 3487 3428 3493
rect 2819 3442 2859 3446
rect 2824 3431 2859 3435
rect 1301 3423 1318 3429
rect 3853 3429 3859 3666
rect 1011 2602 1161 2699
rect 1025 2471 1040 2477
rect 1034 2372 1040 2471
rect 1071 2229 1077 2602
rect 1312 2378 1318 3423
rect 2824 3421 2859 3425
rect 3853 3423 3975 3429
rect 2817 3411 2859 3415
rect 2820 3400 2859 3404
rect 2820 3390 2859 3394
rect 2823 3382 2859 3386
rect 2824 3371 2859 3375
rect 3853 3129 3859 3423
rect 3853 3123 3975 3129
rect 3853 2829 3859 3123
rect 3853 2823 3975 2829
rect 3853 2529 3859 2823
rect 3853 2523 3975 2529
rect 1091 2372 1519 2378
rect 1513 2330 1519 2372
rect 1513 2324 1557 2330
rect 1071 2223 1581 2229
rect 1071 1935 1077 2223
rect 1019 1929 1089 1935
rect 1083 1476 1089 1929
rect 3853 1929 3859 2523
rect 3853 1923 3975 1929
rect 3378 1723 3444 1729
rect 1073 1470 1089 1476
rect 1073 1070 1079 1470
rect 3438 1172 3444 1723
rect 3853 1629 3859 1923
rect 3853 1623 3975 1629
rect 3522 1347 3742 1353
rect 3853 1329 3859 1623
rect 3853 1323 3975 1329
rect 3438 1166 3497 1172
rect 2302 1081 2398 1134
rect 1329 1075 2398 1081
rect 1073 1064 1629 1070
rect 1073 1035 1079 1064
rect 1019 1029 1079 1035
rect 1029 1019 1035 1029
rect 1623 1025 1629 1064
rect 1923 1025 1929 1075
rect 2302 1031 2398 1075
rect 3491 1031 3497 1166
rect 3853 1031 3859 1323
rect 2302 1025 3975 1031
rect 2302 1012 2398 1025
<< m2contact >>
rect 1023 3975 1029 3981
rect 1323 3975 1329 3981
rect 1623 3975 1629 3981
rect 1923 3975 1929 3981
rect 2223 3975 2229 3981
rect 2523 3975 2529 3981
rect 3123 3975 3129 3981
rect 1019 3723 1025 3729
rect 1019 3423 1025 3429
rect 1168 3744 1174 3750
rect 3423 3975 3429 3981
rect 3723 3975 3729 3981
rect 3975 3723 3981 3729
rect 2815 3442 2819 3446
rect 2859 3442 2863 3446
rect 2820 3431 2824 3435
rect 2859 3431 2863 3435
rect 1295 3423 1301 3429
rect 1019 2471 1025 2477
rect 1040 2372 1046 2378
rect 2820 3421 2824 3425
rect 2859 3421 2863 3425
rect 3975 3423 3981 3429
rect 2813 3411 2817 3415
rect 2859 3411 2863 3415
rect 2816 3400 2820 3404
rect 2859 3400 2863 3404
rect 2816 3390 2820 3394
rect 2859 3390 2863 3394
rect 2819 3382 2823 3386
rect 2859 3382 2863 3386
rect 2820 3371 2824 3375
rect 2859 3371 2863 3375
rect 3975 3123 3981 3129
rect 3975 2823 3981 2829
rect 3975 2523 3981 2529
rect 1085 2372 1091 2378
rect 1019 1923 1025 1929
rect 3975 1923 3981 1929
rect 3975 1623 3981 1629
rect 3516 1347 3522 1353
rect 3742 1347 3748 1353
rect 3975 1323 3981 1329
rect 1323 1075 1329 1081
rect 1019 1023 1025 1029
rect 1623 1019 1629 1025
rect 1923 1019 1929 1025
rect 1029 1013 1035 1019
rect 2523 1019 2529 1025
rect 2823 1019 2829 1025
rect 3123 1019 3129 1025
rect 3423 1019 3429 1025
rect 3723 1019 3729 1025
rect 3975 1023 3981 1029
<< metal2 >>
rect 1162 3729 1168 3750
rect 1025 3723 1168 3729
rect 1262 3726 1265 3981
rect 1563 3748 1566 3981
rect 1863 3772 1866 3981
rect 2163 3814 2166 3981
rect 2460 3814 2463 3981
rect 2163 3811 2412 3814
rect 1863 3769 2396 3772
rect 1563 3745 2380 3748
rect 1262 3723 2364 3726
rect 1025 3423 1295 3429
rect 1049 3129 1055 3423
rect 2361 3296 2364 3723
rect 2377 3296 2380 3745
rect 2393 3294 2396 3769
rect 2409 3296 2412 3811
rect 2433 3811 2463 3814
rect 2433 3296 2436 3811
rect 2760 3771 2763 3981
rect 2457 3768 2763 3771
rect 2457 3296 2460 3768
rect 3361 3648 3364 3981
rect 2833 3645 3364 3648
rect 2649 3442 2815 3445
rect 2649 3296 2652 3442
rect 2665 3431 2820 3434
rect 2665 3296 2668 3431
rect 2681 3421 2820 3424
rect 2681 3296 2684 3421
rect 2721 3411 2813 3414
rect 2721 3296 2724 3411
rect 2745 3400 2816 3403
rect 2745 3296 2748 3400
rect 2785 3390 2816 3393
rect 2785 3296 2788 3390
rect 2801 3382 2819 3385
rect 2801 3296 2804 3382
rect 2817 3296 2820 3375
rect 2833 3296 2836 3645
rect 3663 3618 3666 3981
rect 2849 3615 3666 3618
rect 3712 3746 3981 3750
rect 2849 3296 2852 3615
rect 3712 3446 3716 3746
rect 2863 3442 3716 3446
rect 3811 3445 3981 3449
rect 3811 3435 3815 3445
rect 2863 3431 3815 3435
rect 2863 3421 3815 3425
rect 2863 3411 3794 3415
rect 2863 3400 3776 3404
rect 2863 3390 3759 3394
rect 2863 3382 3748 3386
rect 2863 3371 3733 3375
rect 1017 3123 1055 3129
rect 1048 2829 1054 3123
rect 1019 2823 1054 2829
rect 3399 2606 3624 2614
rect 1075 2588 1533 2593
rect 1075 2455 1080 2588
rect 1019 2450 1080 2455
rect 1111 2478 1538 2483
rect 1046 2372 1085 2378
rect 1111 2166 1116 2478
rect 1019 2161 1116 2166
rect 1151 2393 1540 2394
rect 1151 2389 1538 2393
rect 1151 1653 1156 2389
rect 1533 2388 1538 2389
rect 1533 2387 1540 2388
rect 3399 2328 3516 2334
rect 1019 1648 1156 1653
rect 1186 2318 1538 2323
rect 1186 1352 1191 2318
rect 1019 1347 1191 1352
rect 1208 2148 1538 2153
rect 1208 1264 1213 2148
rect 1019 1259 1213 1264
rect 1745 1102 1748 1657
rect 2105 1106 2108 1656
rect 1262 1099 1748 1102
rect 1820 1103 2108 1106
rect 1262 1019 1265 1099
rect 1323 1019 1329 1075
rect 1820 1070 1823 1103
rect 2185 1086 2188 1656
rect 1348 1067 1823 1070
rect 1861 1083 2188 1086
rect 1348 1019 1351 1067
rect 1861 1019 1864 1083
rect 2313 1062 2316 1656
rect 1946 1059 2316 1062
rect 2697 1061 2700 1656
rect 2737 1064 2740 1656
rect 3510 1347 3516 2328
rect 3616 1111 3624 2606
rect 3445 1103 3624 1111
rect 2737 1061 2848 1064
rect 1946 1019 1949 1059
rect 2547 1058 2700 1061
rect 2547 1019 2550 1058
rect 2845 1019 2848 1061
rect 3445 1019 3453 1103
rect 3729 1053 3733 3371
rect 3744 1652 3748 3382
rect 3755 1952 3759 3390
rect 3772 2552 3776 3400
rect 3790 2853 3794 3411
rect 3811 3151 3815 3421
rect 3811 3147 3981 3151
rect 3790 2849 3981 2853
rect 3772 2548 3981 2552
rect 3755 1948 3981 1952
rect 3744 1648 3981 1652
rect 3748 1347 3981 1353
rect 3729 1049 3981 1053
<< m3contact >>
rect 3392 2606 3399 2614
rect 1533 2588 1538 2593
rect 1538 2478 1543 2483
rect 1538 2388 1543 2393
rect 3393 2328 3399 2334
rect 1538 2148 1543 2153
<< metal3 >>
rect 3391 2614 3401 2615
rect 3391 2606 3392 2614
rect 3399 2606 3401 2614
rect 3391 2605 3401 2606
rect 1532 2593 1539 2594
rect 1532 2588 1533 2593
rect 1538 2588 1543 2593
rect 1532 2587 1539 2588
rect 1537 2483 1544 2485
rect 1537 2478 1538 2483
rect 1543 2478 1544 2483
rect 1537 2477 1544 2478
rect 1537 2393 1544 2394
rect 1537 2388 1538 2393
rect 1543 2388 1544 2393
rect 1537 2387 1544 2388
rect 3391 2334 3400 2335
rect 3391 2328 3393 2334
rect 3399 2328 3400 2334
rect 3391 2327 3400 2328
rect 1537 2323 1543 2324
rect 1537 2318 1538 2323
rect 1537 2317 1543 2318
rect 1537 2153 1544 2154
rect 1537 2148 1538 2153
rect 1543 2148 1544 2153
rect 1537 2147 1544 2148
<< rmetal3 >>
rect 1538 2318 1543 2323
use UART  UART_0
timestamp 1554898959
transform 1 0 1543 0 1 1656
box 0 0 1850 1640
use PadFrame  PadFrame_0
timestamp 1554896825
transform 1 0 2500 0 1 2500
box -2500 -2500 2500 2500
<< labels >>
rlabel metal2 2363 3317 2363 3317 1 tx_data[3]
rlabel metal2 2378 3317 2378 3317 1 tx_data[6]
rlabel metal2 2394 3317 2394 3317 1 tx_data[7]
rlabel metal2 2411 3317 2411 3317 1 tx_data[2]
rlabel metal2 2435 3317 2435 3317 1 tx_data[4]
rlabel metal2 2458 3317 2458 3317 1 tx_data[5]
rlabel metal2 2851 3319 2851 3319 1 tx_data[0]
rlabel metal2 2834 3319 2834 3319 1 tx_data[1]
rlabel metal2 2651 3307 2651 3307 1 rxrxout[0]
rlabel metal2 2667 3308 2667 3308 1 rxrxout[6]
rlabel metal2 2683 3308 2683 3308 1 rxrxout[7]
rlabel metal2 1747 1632 1747 1632 1 tx_rdy
rlabel metal2 2107 1632 2107 1632 1 rx_rdy
rlabel metal2 2186 1633 2186 1633 1 reset
rlabel metal2 2699 1623 2699 1623 1 rx_idle
rlabel metal2 2738 1623 2738 1623 1 rx_busy
rlabel metal2 1492 2590 1492 2590 1 tx_idle
rlabel metal2 1494 2480 1494 2480 1 clkb
rlabel metal2 1494 2393 1494 2393 1 tx_error
rlabel metal2 1500 2320 1500 2320 1 tx_busy
rlabel metal2 1514 2151 1514 2151 1 clka
rlabel metal2 2314 1641 2314 1641 1 tx_done
rlabel metal1 1088 2652 1088 2652 1 GND
rlabel metal1 2348 1080 2348 1080 1 VDD
rlabel metal2 1463 2590 1463 2590 1 p_tx_idle
rlabel metal2 1471 2480 1471 2480 1 p_clkb
rlabel metal2 1462 2391 1462 2391 1 p_tx_error
rlabel metal2 1460 2320 1460 2320 1 p_tx_busy
rlabel metal2 1468 2151 1468 2151 1 p_clka
rlabel metal2 1746 1610 1746 1610 1 p_tx_rdy
rlabel metal2 2107 1603 2107 1603 1 p_rx_rdy
rlabel metal2 2186 1605 2186 1605 1 p_reset
rlabel metal2 2314 1605 2314 1605 1 p_tx_done
rlabel metal2 2698 1612 2698 1612 1 p_tx_idle
rlabel metal2 2739 1615 2739 1615 1 p_rx_busy
rlabel metal2 3438 2331 3438 2331 1 p_rx_error
rlabel metal2 3417 2610 3417 2610 1 p_rx_done
rlabel metal2 2850 3305 2850 3305 1 p_tx_data[0]
rlabel metal2 2834 3306 2834 3306 1 p_tx_data[1]
rlabel metal2 2818 3301 2818 3301 1 rxrxout[1]
rlabel metal2 2803 3301 2803 3301 1 rxrxout[2]
rlabel metal2 2786 3302 2786 3302 1 rxrxout[3]
rlabel metal2 2818 3308 2818 3308 1 p_rxrxout[1]
rlabel metal2 2802 3307 2802 3307 1 p_rxrxout[2]
rlabel metal2 2786 3308 2786 3308 1 p_rxrxout[3]
rlabel metal2 2747 3300 2747 3300 1 rxrxout[5]
rlabel metal2 2722 3300 2722 3300 1 rxrxout[4]
rlabel metal2 2747 3307 2747 3307 1 p_rxrxout[5]
rlabel metal2 2722 3309 2722 3309 1 p_rxrxout[4]
rlabel metal2 2682 3320 2682 3320 1 p_rxrxout[7]
rlabel metal2 2666 3318 2666 3318 1 p_rxrxout[6]
rlabel metal2 2651 3317 2651 3317 1 p_rxrxout[0]
rlabel metal2 2458 3310 2458 3310 1 p_tx_data[5]
rlabel metal2 2434 3310 2434 3310 1 p_tx_data[4]
rlabel metal2 2410 3309 2410 3309 1 p_tx_data[2]
rlabel metal2 2395 3309 2395 3309 1 p_tx_data[7]
rlabel metal2 2378 3311 2378 3311 1 p_tx_data[6]
rlabel metal2 2363 3309 2363 3309 1 p_tx_data[3]
<< end >>
