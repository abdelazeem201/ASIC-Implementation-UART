magic
tech scmos
timestamp 1555513135
<< metal1 >>
rect 14 1607 1835 1627
rect 38 1583 1811 1603
rect 38 1567 1811 1573
rect 402 1543 412 1546
rect 354 1526 357 1534
rect 370 1533 420 1536
rect 468 1533 533 1536
rect 564 1533 605 1536
rect 730 1526 733 1534
rect 746 1533 804 1536
rect 818 1533 828 1536
rect 860 1533 901 1536
rect 1036 1533 1053 1536
rect 1154 1533 1172 1536
rect 1276 1533 1293 1536
rect 1420 1533 1437 1536
rect 818 1526 821 1533
rect 1450 1526 1453 1536
rect 252 1523 277 1526
rect 308 1523 357 1526
rect 364 1523 397 1526
rect 436 1523 445 1526
rect 660 1523 685 1526
rect 716 1523 733 1526
rect 740 1523 749 1526
rect 812 1523 821 1526
rect 938 1523 964 1526
rect 468 1513 493 1516
rect 1106 1513 1124 1516
rect 1138 1506 1141 1525
rect 1162 1523 1188 1526
rect 1314 1523 1324 1526
rect 1378 1523 1396 1526
rect 1450 1523 1460 1526
rect 1498 1523 1516 1526
rect 1562 1523 1580 1526
rect 1162 1506 1165 1523
rect 1138 1503 1165 1506
rect 14 1467 1835 1473
rect 1186 1433 1205 1436
rect 300 1423 333 1426
rect 460 1423 533 1426
rect 1202 1425 1205 1433
rect 1498 1416 1501 1425
rect 116 1413 141 1416
rect 196 1413 245 1416
rect 250 1413 284 1416
rect 314 1413 340 1416
rect 522 1413 540 1416
rect 554 1413 564 1416
rect 652 1413 677 1416
rect 778 1413 788 1416
rect 820 1413 837 1416
rect 898 1413 956 1416
rect 988 1413 1021 1416
rect 1050 1413 1077 1416
rect 1154 1413 1172 1416
rect 1484 1413 1501 1416
rect 1530 1413 1564 1416
rect 674 1406 677 1413
rect 162 1403 172 1406
rect 204 1403 276 1406
rect 348 1403 365 1406
rect 378 1403 428 1406
rect 458 1403 532 1406
rect 546 1403 556 1406
rect 602 1403 644 1406
rect 674 1403 684 1406
rect 716 1403 749 1406
rect 906 1403 948 1406
rect 1074 1405 1077 1413
rect 1124 1403 1133 1406
rect 1140 1403 1165 1406
rect 1458 1403 1476 1406
rect 1692 1403 1701 1406
rect 1162 1393 1165 1403
rect 38 1367 1811 1373
rect 394 1343 436 1346
rect 1028 1343 1037 1346
rect 242 1333 252 1336
rect 314 1333 332 1336
rect 444 1333 469 1336
rect 514 1333 532 1336
rect 556 1333 605 1336
rect 260 1323 285 1326
rect 290 1323 324 1326
rect 356 1323 365 1326
rect 522 1323 540 1326
rect 642 1323 645 1334
rect 650 1333 660 1336
rect 698 1333 740 1336
rect 762 1333 772 1336
rect 908 1333 925 1336
rect 930 1333 940 1336
rect 988 1333 1005 1336
rect 1020 1333 1053 1336
rect 1202 1333 1236 1336
rect 1442 1333 1492 1336
rect 1626 1333 1644 1336
rect 1658 1333 1668 1336
rect 658 1323 668 1326
rect 722 1323 732 1326
rect 780 1323 789 1326
rect 858 1323 884 1326
rect 964 1323 1012 1326
rect 1218 1323 1221 1333
rect 1330 1323 1380 1326
rect 1410 1323 1420 1326
rect 1482 1323 1500 1326
rect 1506 1323 1532 1326
rect 1562 1323 1588 1326
rect 1652 1323 1669 1326
rect 1684 1323 1717 1326
rect 290 1316 293 1323
rect 1482 1316 1485 1323
rect 138 1313 164 1316
rect 188 1313 197 1316
rect 268 1313 293 1316
rect 556 1313 589 1316
rect 1436 1313 1485 1316
rect 1666 1315 1669 1323
rect 836 1303 853 1306
rect 14 1267 1835 1273
rect 284 1223 316 1226
rect 418 1216 421 1225
rect 1674 1216 1677 1225
rect 170 1213 180 1216
rect 194 1213 212 1216
rect 244 1213 253 1216
rect 266 1213 276 1216
rect 330 1213 405 1216
rect 418 1213 428 1216
rect 434 1213 444 1216
rect 476 1213 517 1216
rect 524 1213 548 1216
rect 562 1213 580 1216
rect 610 1213 628 1216
rect 634 1213 652 1216
rect 724 1213 773 1216
rect 890 1213 964 1216
rect 1194 1213 1212 1216
rect 1266 1213 1284 1216
rect 1452 1213 1477 1216
rect 1514 1213 1524 1216
rect 1530 1213 1548 1216
rect 1660 1213 1677 1216
rect 1692 1213 1733 1216
rect 218 1203 236 1206
rect 250 1203 268 1206
rect 402 1205 405 1213
rect 436 1203 445 1206
rect 474 1203 516 1206
rect 660 1203 693 1206
rect 786 1203 796 1206
rect 828 1203 860 1206
rect 908 1203 917 1206
rect 930 1203 956 1206
rect 980 1203 997 1206
rect 1116 1203 1165 1206
rect 1396 1203 1413 1206
rect 1642 1203 1652 1206
rect 38 1167 1811 1173
rect 282 1143 324 1146
rect 1442 1143 1469 1146
rect 1466 1136 1469 1143
rect 108 1133 125 1136
rect 170 1133 220 1136
rect 244 1135 301 1136
rect 242 1133 301 1135
rect 340 1133 349 1136
rect 564 1133 573 1136
rect 900 1133 933 1136
rect 116 1123 157 1126
rect 164 1123 181 1126
rect 242 1123 245 1133
rect 1186 1126 1189 1135
rect 1218 1133 1236 1136
rect 1354 1126 1357 1135
rect 1436 1133 1461 1136
rect 1466 1133 1476 1136
rect 1490 1126 1493 1135
rect 1666 1126 1669 1135
rect 290 1123 324 1126
rect 676 1123 701 1126
rect 810 1123 820 1126
rect 954 1123 964 1126
rect 994 1123 1020 1126
rect 1092 1123 1117 1126
rect 1148 1123 1189 1126
rect 1234 1123 1244 1126
rect 1292 1123 1317 1126
rect 1348 1123 1357 1126
rect 1402 1123 1477 1126
rect 1484 1123 1493 1126
rect 1604 1123 1629 1126
rect 1660 1123 1669 1126
rect 1714 1126 1717 1135
rect 1722 1133 1740 1136
rect 1714 1123 1748 1126
rect 564 1113 597 1116
rect 914 1113 940 1116
rect 1372 1113 1397 1116
rect 14 1067 1835 1073
rect 116 1033 125 1036
rect 132 1023 157 1026
rect 892 1023 917 1026
rect 970 1016 973 1025
rect 1146 1023 1156 1026
rect 1356 1023 1365 1026
rect 244 1013 285 1016
rect 330 1013 340 1016
rect 700 1013 709 1016
rect 812 1013 821 1016
rect 874 1013 884 1016
rect 922 1013 956 1016
rect 970 1013 988 1016
rect 994 1013 1020 1016
rect 1050 1013 1076 1016
rect 1124 1013 1157 1016
rect 1164 1013 1173 1016
rect 1250 1013 1276 1016
rect 1314 1013 1340 1016
rect 1404 1013 1429 1016
rect 1460 1013 1477 1016
rect 1612 1013 1637 1016
rect 1668 1013 1677 1016
rect 1684 1013 1709 1016
rect 138 1003 172 1006
rect 194 1003 236 1006
rect 274 1003 292 1006
rect 356 1003 389 1006
rect 572 1003 605 1006
rect 890 1003 948 1006
rect 972 1003 981 1006
rect 994 1005 997 1013
rect 1204 1003 1213 1006
rect 1322 1003 1332 1006
rect 1482 1003 1500 1006
rect 1674 1005 1677 1013
rect 1698 1003 1716 1006
rect 1748 1003 1757 1006
rect 138 993 164 996
rect 38 967 1811 973
rect 322 926 325 934
rect 338 933 404 936
rect 434 926 437 934
rect 452 933 485 936
rect 618 926 621 934
rect 682 933 700 936
rect 724 933 733 936
rect 786 926 789 934
rect 794 933 844 936
rect 892 933 933 936
rect 986 933 1004 936
rect 1066 933 1092 936
rect 1236 933 1245 936
rect 1466 926 1469 945
rect 66 923 76 926
rect 170 923 188 926
rect 210 923 325 926
rect 332 923 357 926
rect 434 923 453 926
rect 612 923 621 926
rect 722 923 748 926
rect 762 923 780 926
rect 786 923 813 926
rect 834 923 852 926
rect 866 923 884 926
rect 980 923 997 926
rect 1060 923 1093 926
rect 1148 923 1173 926
rect 1210 923 1220 926
rect 1234 923 1252 926
rect 1404 923 1413 926
rect 1436 923 1469 926
rect 1506 923 1540 926
rect 1570 923 1573 934
rect 1620 933 1629 936
rect 1650 926 1653 934
rect 1722 933 1748 936
rect 1644 923 1653 926
rect 210 916 213 923
rect 196 913 213 916
rect 340 913 381 916
rect 762 915 765 923
rect 866 915 869 923
rect 1236 913 1245 916
rect 14 867 1835 873
rect 316 833 325 836
rect 330 833 349 836
rect 260 823 308 826
rect 330 825 333 833
rect 364 823 405 826
rect 508 823 541 826
rect 1146 823 1180 826
rect 1474 823 1492 826
rect 538 816 541 823
rect 130 813 173 816
rect 132 803 141 806
rect 170 805 173 813
rect 194 805 197 816
rect 202 813 252 816
rect 450 813 492 816
rect 538 813 556 816
rect 924 813 933 816
rect 980 813 1013 816
rect 1044 813 1069 816
rect 1124 813 1181 816
rect 1196 813 1213 816
rect 1308 813 1333 816
rect 1388 813 1421 816
rect 1444 813 1485 816
rect 1540 813 1549 816
rect 1572 813 1597 816
rect 1418 806 1421 813
rect 1634 806 1637 816
rect 1644 813 1653 816
rect 226 803 244 806
rect 474 803 484 806
rect 508 803 541 806
rect 946 803 956 806
rect 986 803 1020 806
rect 1170 803 1180 806
rect 1204 803 1213 806
rect 1410 805 1421 806
rect 1410 803 1420 805
rect 1538 803 1548 806
rect 1596 805 1637 806
rect 1674 805 1677 816
rect 1716 813 1733 816
rect 1596 803 1636 805
rect 38 767 1811 773
rect 282 726 285 734
rect 122 723 148 726
rect 276 723 285 726
rect 292 723 317 726
rect 426 716 429 734
rect 482 726 485 734
rect 498 733 532 736
rect 564 733 573 736
rect 706 726 709 734
rect 714 733 732 736
rect 794 733 804 736
rect 828 733 853 736
rect 954 733 964 736
rect 994 733 1028 736
rect 1058 733 1084 736
rect 1458 733 1468 736
rect 436 723 485 726
rect 498 723 540 726
rect 612 723 637 726
rect 706 723 812 726
rect 988 723 1021 726
rect 1052 723 1085 726
rect 1092 723 1109 726
rect 1196 723 1213 726
rect 1218 723 1244 726
rect 1364 723 1373 726
rect 1452 723 1469 726
rect 1490 723 1493 734
rect 1522 733 1548 736
rect 1660 733 1668 736
rect 1514 723 1540 726
rect 1588 723 1645 726
rect 1652 723 1669 726
rect 1676 723 1701 726
rect 1716 723 1733 726
rect 1754 723 1757 734
rect 348 713 429 716
rect 828 713 853 716
rect 1100 713 1133 716
rect 1594 713 1644 716
rect 1690 713 1700 716
rect 330 703 340 706
rect 850 703 853 713
rect 14 667 1835 673
rect 356 623 405 626
rect 506 623 524 626
rect 978 623 1012 626
rect 170 613 188 616
rect 306 613 324 616
rect 482 613 492 616
rect 540 613 564 616
rect 722 613 740 616
rect 804 613 813 616
rect 820 613 837 616
rect 850 613 900 616
rect 948 613 957 616
rect 964 613 973 616
rect 1010 613 1020 616
rect 1050 613 1149 616
rect 1146 606 1149 613
rect 1218 606 1221 616
rect 1282 613 1308 616
rect 1490 613 1500 616
rect 1572 613 1597 616
rect 1594 606 1597 613
rect 1674 613 1733 616
rect 1740 613 1757 616
rect 1674 606 1677 613
rect 282 603 316 606
rect 442 603 468 606
rect 580 603 621 606
rect 754 603 796 606
rect 852 603 869 606
rect 908 603 933 606
rect 1146 603 1172 606
rect 1204 603 1221 606
rect 1404 603 1429 606
rect 1474 603 1492 606
rect 1554 603 1564 606
rect 1594 603 1636 606
rect 1652 603 1677 606
rect 1682 603 1692 606
rect 1730 605 1733 613
rect 442 595 445 603
rect 38 567 1811 573
rect 138 533 165 536
rect 356 533 381 536
rect 450 533 468 536
rect 612 533 628 536
rect 900 533 940 536
rect 1028 533 1044 536
rect 74 523 92 526
rect 138 525 141 533
rect 1306 526 1309 535
rect 1386 533 1436 536
rect 1468 533 1493 536
rect 1522 533 1556 536
rect 1580 533 1636 536
rect 1666 533 1692 536
rect 1714 526 1717 535
rect 146 523 172 526
rect 290 523 316 526
rect 354 523 429 526
rect 522 523 548 526
rect 594 523 604 526
rect 644 523 669 526
rect 708 523 717 526
rect 764 523 773 526
rect 874 523 884 526
rect 906 523 948 526
rect 954 523 1020 526
rect 1122 523 1132 526
rect 1244 523 1269 526
rect 1300 523 1309 526
rect 1380 523 1405 526
rect 1418 523 1453 526
rect 1460 523 1469 526
rect 1516 523 1557 526
rect 1572 523 1629 526
rect 1634 523 1644 526
rect 1714 523 1725 526
rect 1738 523 1748 526
rect 452 513 469 516
rect 1388 513 1397 516
rect 1450 515 1453 523
rect 1530 513 1556 516
rect 14 467 1835 473
rect 116 433 133 436
rect 978 433 1020 436
rect 1098 433 1132 436
rect 98 423 108 426
rect 132 423 149 426
rect 978 423 1004 426
rect 1098 423 1116 426
rect 1162 423 1228 426
rect 1314 423 1340 426
rect 1314 416 1317 423
rect 1506 416 1509 425
rect 204 413 221 416
rect 322 413 332 416
rect 362 413 404 416
rect 460 413 469 416
rect 506 413 532 416
rect 612 413 621 416
rect 668 413 701 416
rect 954 413 972 416
rect 1034 413 1084 416
rect 1236 413 1253 416
rect 1284 413 1317 416
rect 1356 413 1436 416
rect 1506 413 1516 416
rect 1628 413 1645 416
rect 1652 413 1677 416
rect 1716 413 1725 416
rect 234 403 244 406
rect 306 403 324 406
rect 356 403 373 406
rect 426 403 436 406
rect 860 403 901 406
rect 932 403 949 406
rect 1250 403 1260 406
rect 1292 403 1317 406
rect 1330 403 1340 406
rect 1364 403 1429 406
rect 1458 403 1492 406
rect 1460 393 1485 396
rect 38 367 1811 373
rect 602 343 636 346
rect 1524 343 1541 346
rect 1538 336 1541 343
rect 306 333 324 336
rect 618 333 644 336
rect 714 333 725 336
rect 1146 333 1164 336
rect 1212 333 1245 336
rect 1250 333 1276 336
rect 1460 333 1477 336
rect 1490 333 1508 336
rect 1538 333 1564 336
rect 1594 333 1644 336
rect 290 323 332 326
rect 378 323 404 326
rect 596 323 637 326
rect 652 323 661 326
rect 714 325 717 333
rect 1172 323 1189 326
rect 1290 323 1356 326
rect 1394 323 1428 326
rect 1442 323 1452 326
rect 122 313 173 316
rect 210 313 244 316
rect 722 313 804 316
rect 818 313 828 316
rect 1044 313 1069 316
rect 1100 313 1133 316
rect 1186 315 1189 323
rect 1594 315 1597 333
rect 90 303 180 306
rect 252 303 269 306
rect 1050 303 1092 306
rect 14 267 1835 273
rect 1058 233 1092 236
rect 1356 233 1381 236
rect 652 223 685 226
rect 716 223 804 226
rect 1050 223 1076 226
rect 1100 223 1133 226
rect 1308 223 1348 226
rect 1362 223 1372 226
rect 1394 223 1444 226
rect 1468 223 1493 226
rect 1524 223 1549 226
rect 124 213 165 216
rect 170 213 212 216
rect 372 213 437 216
rect 644 213 661 216
rect 940 213 957 216
rect 1186 213 1204 216
rect 1242 213 1292 216
rect 1530 213 1572 216
rect 1578 213 1645 216
rect 1772 213 1781 216
rect 74 203 108 206
rect 234 203 252 206
rect 444 203 461 206
rect 548 203 629 206
rect 954 203 1012 206
rect 1482 203 1500 206
rect 1524 203 1541 206
rect 1578 205 1581 213
rect 1586 203 1620 206
rect 394 193 436 196
rect 38 167 1811 173
rect 1164 143 1189 146
rect 1186 136 1189 143
rect 172 133 181 136
rect 258 133 332 136
rect 356 133 381 136
rect 580 133 589 136
rect 684 133 701 136
rect 738 133 748 136
rect 802 133 812 136
rect 970 133 980 136
rect 1122 133 1156 136
rect 1186 133 1196 136
rect 1386 133 1436 136
rect 1666 126 1669 136
rect 330 123 340 126
rect 492 123 549 126
rect 676 123 797 126
rect 988 123 1021 126
rect 1116 123 1148 126
rect 1210 123 1228 126
rect 1388 123 1397 126
rect 1466 123 1516 126
rect 1570 123 1596 126
rect 1644 123 1669 126
rect 236 113 325 116
rect 178 103 228 106
rect 202 93 205 103
rect 14 67 1835 73
rect 38 37 1811 57
rect 14 13 1835 33
<< metal2 >>
rect 14 13 34 1627
rect 38 37 58 1603
rect 362 1576 365 1640
rect 354 1573 365 1576
rect 162 1533 165 1546
rect 82 1493 85 1526
rect 138 1513 141 1526
rect 106 1403 109 1426
rect 138 1313 141 1416
rect 162 1383 165 1496
rect 178 1413 181 1426
rect 186 1403 189 1516
rect 202 1496 205 1546
rect 226 1533 229 1546
rect 354 1536 357 1573
rect 410 1556 413 1640
rect 410 1553 421 1556
rect 354 1533 373 1536
rect 274 1513 277 1526
rect 202 1493 213 1496
rect 210 1426 213 1493
rect 202 1423 213 1426
rect 74 1143 77 1216
rect 130 1193 133 1216
rect 154 1146 157 1366
rect 202 1363 205 1423
rect 170 1213 173 1326
rect 178 1293 181 1306
rect 194 1223 197 1316
rect 226 1296 229 1406
rect 242 1403 245 1416
rect 242 1313 245 1336
rect 178 1213 197 1216
rect 98 1143 109 1146
rect 122 1116 125 1136
rect 138 1126 141 1146
rect 114 1113 125 1116
rect 134 1123 141 1126
rect 146 1143 157 1146
rect 170 1146 173 1206
rect 194 1193 197 1206
rect 170 1143 181 1146
rect 202 1143 205 1206
rect 218 1203 221 1296
rect 226 1293 237 1296
rect 234 1226 237 1293
rect 226 1223 237 1226
rect 226 1193 229 1223
rect 250 1213 253 1416
rect 266 1213 269 1426
rect 274 1403 293 1406
rect 298 1403 301 1516
rect 314 1403 317 1416
rect 330 1406 333 1426
rect 330 1403 341 1406
rect 290 1386 293 1403
rect 290 1383 301 1386
rect 282 1323 285 1366
rect 298 1316 301 1383
rect 290 1313 301 1316
rect 114 1056 117 1113
rect 114 1053 125 1056
rect 122 1033 125 1053
rect 134 1026 137 1123
rect 106 966 109 1026
rect 134 1023 141 1026
rect 122 996 125 1016
rect 138 1003 141 1023
rect 146 1006 149 1143
rect 154 1133 173 1136
rect 154 1113 157 1126
rect 178 1123 181 1143
rect 210 1116 213 1136
rect 202 1113 213 1116
rect 202 1056 205 1113
rect 218 1103 221 1116
rect 234 1113 237 1206
rect 250 1136 253 1206
rect 282 1156 285 1226
rect 274 1153 285 1156
rect 250 1133 261 1136
rect 242 1096 245 1126
rect 226 1093 245 1096
rect 154 1013 157 1026
rect 146 1003 157 1006
rect 122 993 141 996
rect 106 963 117 966
rect 66 923 69 936
rect 114 886 117 963
rect 106 883 117 886
rect 66 823 69 866
rect 74 716 77 736
rect 82 723 85 826
rect 106 823 109 883
rect 122 813 125 826
rect 130 813 133 926
rect 154 816 157 1003
rect 162 993 165 1056
rect 202 1053 213 1056
rect 186 1013 189 1036
rect 194 1003 197 1016
rect 178 933 189 936
rect 170 823 173 926
rect 210 923 213 1053
rect 154 813 173 816
rect 186 813 189 836
rect 194 813 197 916
rect 106 803 125 806
rect 90 716 93 726
rect 122 723 125 803
rect 138 793 141 806
rect 170 723 173 813
rect 202 793 205 816
rect 226 803 229 1093
rect 258 1086 261 1133
rect 250 1083 261 1086
rect 250 1013 253 1083
rect 274 1003 277 1153
rect 282 1133 285 1146
rect 290 1103 293 1313
rect 314 1193 317 1336
rect 322 1286 325 1326
rect 338 1323 341 1403
rect 354 1393 357 1533
rect 394 1506 397 1526
rect 386 1503 397 1506
rect 386 1426 389 1503
rect 402 1436 405 1546
rect 402 1433 409 1436
rect 386 1423 397 1426
rect 346 1333 349 1346
rect 362 1323 365 1406
rect 378 1383 381 1406
rect 394 1343 397 1423
rect 406 1386 409 1433
rect 418 1403 421 1553
rect 434 1533 445 1536
rect 530 1533 533 1546
rect 442 1513 445 1526
rect 434 1403 437 1416
rect 450 1413 453 1526
rect 490 1503 493 1516
rect 514 1436 517 1516
rect 538 1513 541 1536
rect 546 1533 549 1640
rect 730 1556 733 1576
rect 546 1446 549 1526
rect 562 1503 565 1516
rect 546 1443 557 1446
rect 506 1433 517 1436
rect 402 1383 409 1386
rect 402 1363 405 1383
rect 322 1283 333 1286
rect 298 1133 301 1186
rect 282 1013 301 1016
rect 306 1003 309 1116
rect 322 1053 325 1216
rect 330 1213 333 1283
rect 330 1193 333 1206
rect 338 1183 341 1206
rect 338 1156 341 1176
rect 334 1153 341 1156
rect 334 1056 337 1153
rect 346 1133 349 1216
rect 410 1183 413 1216
rect 418 1173 421 1216
rect 434 1213 437 1346
rect 442 1333 445 1406
rect 450 1403 461 1406
rect 450 1323 453 1403
rect 466 1306 469 1336
rect 458 1303 469 1306
rect 458 1236 461 1303
rect 474 1286 477 1426
rect 506 1356 509 1433
rect 530 1423 549 1426
rect 506 1353 517 1356
rect 514 1333 517 1353
rect 522 1323 525 1416
rect 554 1413 557 1443
rect 530 1403 549 1406
rect 530 1333 541 1336
rect 546 1333 549 1403
rect 474 1283 485 1286
rect 458 1233 469 1236
rect 442 1196 445 1206
rect 450 1203 453 1216
rect 458 1196 461 1216
rect 442 1193 461 1196
rect 466 1193 469 1233
rect 482 1226 485 1283
rect 474 1223 485 1226
rect 474 1186 477 1223
rect 514 1213 517 1226
rect 530 1223 533 1236
rect 474 1183 481 1186
rect 334 1053 341 1056
rect 250 813 253 946
rect 314 943 317 1016
rect 322 1003 325 1046
rect 330 1013 333 1036
rect 338 1006 341 1053
rect 346 1043 349 1126
rect 410 1056 413 1136
rect 434 1113 437 1126
rect 478 1116 481 1183
rect 490 1123 493 1156
rect 538 1133 541 1333
rect 554 1226 557 1316
rect 554 1223 565 1226
rect 546 1213 565 1216
rect 546 1123 549 1213
rect 562 1193 565 1206
rect 554 1116 557 1186
rect 570 1153 573 1536
rect 586 1313 589 1506
rect 602 1496 605 1536
rect 634 1533 637 1556
rect 722 1553 733 1556
rect 754 1556 757 1626
rect 818 1573 821 1640
rect 754 1553 773 1556
rect 682 1506 685 1526
rect 674 1503 685 1506
rect 602 1493 613 1496
rect 610 1446 613 1493
rect 602 1443 613 1446
rect 602 1403 605 1443
rect 674 1426 677 1503
rect 722 1466 725 1553
rect 746 1533 749 1546
rect 722 1463 733 1466
rect 674 1423 685 1426
rect 682 1406 685 1423
rect 690 1413 693 1456
rect 730 1426 733 1463
rect 706 1413 709 1426
rect 722 1423 733 1426
rect 602 1333 605 1346
rect 586 1223 589 1236
rect 474 1113 481 1116
rect 538 1113 557 1116
rect 474 1093 477 1113
rect 402 1053 413 1056
rect 330 1003 341 1006
rect 338 923 341 936
rect 354 913 357 1026
rect 386 933 389 1006
rect 402 993 405 1053
rect 538 1046 541 1113
rect 570 1106 573 1136
rect 562 1103 573 1106
rect 538 1043 549 1046
rect 426 996 429 1016
rect 418 993 429 996
rect 338 836 341 846
rect 258 823 261 836
rect 314 833 341 836
rect 290 773 293 826
rect 314 816 317 833
rect 306 813 317 816
rect 74 713 93 716
rect 90 663 93 713
rect 74 286 77 526
rect 82 493 85 616
rect 106 536 109 616
rect 114 543 117 556
rect 122 543 125 666
rect 162 613 165 626
rect 170 536 173 616
rect 194 573 197 736
rect 218 656 221 726
rect 218 653 229 656
rect 226 576 229 653
rect 242 603 245 616
rect 218 573 229 576
rect 98 423 101 536
rect 106 533 117 536
rect 114 523 117 533
rect 130 506 133 536
rect 162 533 173 536
rect 202 536 205 556
rect 202 533 209 536
rect 122 503 133 506
rect 122 456 125 503
rect 122 453 133 456
rect 130 433 133 453
rect 90 303 93 376
rect 74 283 85 286
rect 82 226 85 283
rect 74 223 85 226
rect 74 203 77 223
rect 106 113 109 326
rect 122 313 125 416
rect 130 413 133 426
rect 146 423 149 526
rect 162 516 165 533
rect 162 513 173 516
rect 170 436 173 513
rect 206 486 209 533
rect 162 433 173 436
rect 202 483 209 486
rect 162 373 165 433
rect 178 403 181 416
rect 162 323 173 326
rect 130 203 133 306
rect 162 123 165 216
rect 170 213 173 316
rect 186 313 189 406
rect 202 393 205 483
rect 218 413 221 573
rect 266 566 269 726
rect 274 713 277 726
rect 282 603 285 626
rect 250 563 269 566
rect 250 533 253 563
rect 226 513 229 526
rect 290 523 293 726
rect 306 546 309 813
rect 322 736 325 826
rect 338 823 341 833
rect 314 733 325 736
rect 314 723 317 733
rect 346 726 349 836
rect 354 833 373 836
rect 370 816 373 833
rect 362 813 373 816
rect 362 746 365 813
rect 378 756 381 916
rect 402 896 405 936
rect 410 923 413 936
rect 418 933 421 993
rect 482 933 485 1016
rect 522 1003 525 1026
rect 530 1013 541 1016
rect 546 1013 549 1043
rect 562 1013 565 1103
rect 538 1003 541 1013
rect 426 913 429 926
rect 402 893 413 896
rect 402 763 405 826
rect 410 823 413 893
rect 378 753 389 756
rect 362 743 373 746
rect 330 723 357 726
rect 322 623 325 716
rect 330 703 333 716
rect 354 666 357 723
rect 370 713 373 743
rect 386 706 389 753
rect 418 726 421 836
rect 426 813 429 826
rect 434 823 437 846
rect 450 813 453 926
rect 530 836 533 946
rect 554 923 557 1006
rect 578 966 581 1116
rect 594 1113 597 1246
rect 610 1233 613 1396
rect 618 1323 621 1406
rect 682 1403 701 1406
rect 610 1133 613 1216
rect 626 1213 629 1336
rect 634 1323 637 1336
rect 650 1333 653 1366
rect 642 1313 645 1326
rect 658 1303 661 1326
rect 698 1316 701 1366
rect 722 1346 725 1423
rect 722 1343 733 1346
rect 690 1313 701 1316
rect 690 1246 693 1313
rect 722 1306 725 1326
rect 730 1323 733 1343
rect 690 1243 701 1246
rect 634 1213 637 1226
rect 690 1213 693 1226
rect 570 963 581 966
rect 602 963 605 1126
rect 618 1123 621 1186
rect 626 1066 629 1136
rect 634 1123 637 1206
rect 690 1196 693 1206
rect 698 1203 701 1243
rect 706 1196 709 1216
rect 714 1203 717 1306
rect 722 1303 729 1306
rect 726 1206 729 1303
rect 722 1203 729 1206
rect 690 1193 709 1196
rect 642 1133 645 1146
rect 650 1123 653 1136
rect 698 1133 701 1186
rect 722 1183 725 1203
rect 738 1193 741 1456
rect 746 1403 749 1526
rect 770 1436 773 1553
rect 818 1546 821 1566
rect 814 1543 821 1546
rect 802 1513 805 1536
rect 754 1433 773 1436
rect 746 1313 749 1326
rect 698 1096 701 1126
rect 690 1093 701 1096
rect 626 1063 645 1066
rect 642 1013 645 1063
rect 690 1026 693 1093
rect 706 1033 709 1146
rect 754 1133 757 1433
rect 814 1426 817 1543
rect 834 1536 837 1640
rect 850 1563 853 1640
rect 866 1623 869 1640
rect 890 1623 893 1640
rect 826 1533 837 1536
rect 842 1533 845 1546
rect 814 1423 821 1426
rect 762 1333 765 1346
rect 762 1303 765 1326
rect 770 1213 773 1336
rect 778 1303 781 1416
rect 794 1383 797 1406
rect 802 1403 805 1416
rect 810 1363 813 1406
rect 818 1356 821 1423
rect 802 1353 821 1356
rect 786 1203 789 1326
rect 802 1246 805 1353
rect 818 1326 821 1346
rect 826 1333 829 1533
rect 834 1453 837 1526
rect 850 1513 853 1526
rect 898 1516 901 1536
rect 890 1513 901 1516
rect 890 1456 893 1513
rect 890 1453 901 1456
rect 834 1393 837 1416
rect 814 1323 821 1326
rect 814 1266 817 1323
rect 814 1263 821 1266
rect 802 1243 813 1246
rect 810 1223 813 1243
rect 802 1193 805 1216
rect 818 1213 821 1263
rect 730 1096 733 1126
rect 762 1123 765 1146
rect 722 1093 733 1096
rect 690 1023 701 1026
rect 698 1006 701 1023
rect 706 1013 709 1026
rect 722 1023 725 1093
rect 570 886 573 963
rect 618 943 621 1006
rect 698 1003 709 1006
rect 626 913 629 966
rect 682 916 685 936
rect 714 923 717 1016
rect 730 1003 733 1026
rect 738 1013 741 1036
rect 730 933 733 996
rect 770 993 773 1156
rect 810 1123 813 1206
rect 826 1153 829 1316
rect 834 1233 837 1356
rect 842 1323 845 1436
rect 850 1353 853 1416
rect 874 1413 877 1436
rect 898 1413 901 1453
rect 898 1393 901 1406
rect 906 1403 909 1526
rect 914 1393 917 1640
rect 930 1566 933 1640
rect 922 1563 933 1566
rect 922 1476 925 1563
rect 938 1523 941 1546
rect 922 1473 929 1476
rect 926 1426 929 1473
rect 926 1423 933 1426
rect 858 1336 861 1346
rect 850 1333 861 1336
rect 850 1323 861 1326
rect 850 1313 853 1323
rect 850 1293 853 1306
rect 882 1213 885 1296
rect 890 1213 893 1236
rect 858 1156 861 1206
rect 858 1153 869 1156
rect 818 1013 821 1126
rect 842 1103 845 1136
rect 858 1133 861 1146
rect 866 1123 869 1153
rect 874 1123 877 1136
rect 890 1123 893 1136
rect 906 1126 909 1356
rect 914 1203 917 1386
rect 922 1316 925 1416
rect 930 1363 933 1423
rect 930 1333 933 1346
rect 922 1313 929 1316
rect 926 1226 929 1313
rect 922 1223 929 1226
rect 902 1123 909 1126
rect 786 983 789 1006
rect 738 933 741 946
rect 762 926 765 936
rect 674 913 685 916
rect 570 883 581 886
rect 522 833 533 836
rect 378 703 389 706
rect 402 723 421 726
rect 354 663 365 666
rect 338 633 341 646
rect 330 613 333 626
rect 346 613 349 626
rect 362 606 365 663
rect 298 543 309 546
rect 298 516 301 543
rect 282 513 301 516
rect 210 313 213 406
rect 234 403 237 416
rect 250 323 253 416
rect 218 136 221 206
rect 234 203 237 216
rect 258 213 261 486
rect 282 436 285 513
rect 282 433 293 436
rect 266 396 269 416
rect 266 393 277 396
rect 274 336 277 393
rect 266 333 277 336
rect 266 313 269 333
rect 290 323 293 433
rect 306 333 309 536
rect 322 533 325 606
rect 346 603 365 606
rect 338 533 341 546
rect 330 483 333 526
rect 322 413 325 476
rect 338 403 341 516
rect 346 473 349 603
rect 370 586 373 626
rect 378 613 381 703
rect 402 623 405 723
rect 410 603 413 716
rect 442 703 445 776
rect 474 706 477 806
rect 522 776 525 833
rect 538 803 541 826
rect 546 783 549 806
rect 522 773 533 776
rect 466 703 477 706
rect 466 646 469 703
rect 418 603 421 616
rect 426 613 429 646
rect 466 643 477 646
rect 474 613 477 643
rect 482 623 485 726
rect 362 583 373 586
rect 362 533 365 583
rect 354 493 357 526
rect 346 393 349 416
rect 362 413 365 436
rect 266 196 269 306
rect 338 266 341 336
rect 354 333 357 406
rect 370 403 373 546
rect 378 516 381 536
rect 418 533 421 546
rect 434 533 437 606
rect 442 593 445 606
rect 378 513 389 516
rect 386 436 389 513
rect 378 433 389 436
rect 346 303 349 326
rect 378 323 381 433
rect 322 263 341 266
rect 322 213 325 263
rect 346 203 349 226
rect 362 223 365 236
rect 178 103 181 136
rect 210 133 221 136
rect 258 193 269 196
rect 210 113 213 133
rect 218 113 221 126
rect 202 0 205 96
rect 258 0 261 193
rect 378 133 381 206
rect 394 193 397 416
rect 418 393 421 406
rect 426 403 429 526
rect 442 523 445 546
rect 450 503 453 536
rect 466 513 469 526
rect 474 523 477 536
rect 482 523 485 616
rect 490 556 493 746
rect 498 733 501 766
rect 530 753 533 773
rect 562 743 565 846
rect 578 806 581 883
rect 674 836 677 913
rect 674 833 685 836
rect 618 813 621 826
rect 570 803 581 806
rect 498 706 501 726
rect 538 713 541 726
rect 498 703 509 706
rect 546 703 549 716
rect 506 646 509 703
rect 498 643 509 646
rect 498 603 501 643
rect 490 553 501 556
rect 482 496 485 516
rect 490 503 493 526
rect 498 496 501 553
rect 506 533 509 626
rect 522 523 525 606
rect 546 603 549 626
rect 554 603 557 726
rect 570 703 573 803
rect 586 733 589 776
rect 594 766 597 806
rect 674 783 677 816
rect 594 763 621 766
rect 618 696 621 763
rect 634 723 637 746
rect 666 723 669 736
rect 674 733 677 766
rect 682 723 685 833
rect 690 733 693 746
rect 698 713 701 916
rect 722 913 725 926
rect 754 923 765 926
rect 754 813 757 923
rect 770 843 773 916
rect 794 856 797 946
rect 810 906 813 926
rect 834 923 837 1036
rect 866 1006 869 1016
rect 874 1013 877 1116
rect 902 1046 905 1123
rect 902 1043 909 1046
rect 866 1003 877 1006
rect 874 993 877 1003
rect 890 943 893 1006
rect 866 926 869 936
rect 858 923 869 926
rect 858 906 861 923
rect 810 903 821 906
rect 858 903 869 906
rect 874 903 877 916
rect 794 853 801 856
rect 730 773 733 806
rect 798 776 801 853
rect 818 846 821 903
rect 810 843 821 846
rect 810 793 813 843
rect 866 813 869 903
rect 898 856 901 1026
rect 906 933 909 1043
rect 914 1023 917 1116
rect 922 1013 925 1223
rect 930 1106 933 1206
rect 938 1183 941 1516
rect 946 1353 949 1640
rect 954 1373 957 1546
rect 962 1383 965 1626
rect 970 1543 973 1640
rect 1010 1566 1013 1586
rect 1006 1563 1013 1566
rect 986 1413 989 1536
rect 1006 1506 1009 1563
rect 1018 1513 1021 1640
rect 1090 1623 1093 1640
rect 1006 1503 1013 1506
rect 1010 1403 1013 1503
rect 1026 1436 1029 1546
rect 1018 1433 1029 1436
rect 1018 1413 1021 1433
rect 1042 1413 1045 1526
rect 1050 1523 1053 1536
rect 1050 1413 1053 1446
rect 1018 1393 1021 1406
rect 1066 1403 1069 1566
rect 1090 1413 1093 1606
rect 1106 1543 1109 1640
rect 1122 1603 1125 1640
rect 1138 1536 1141 1640
rect 1162 1626 1165 1640
rect 1154 1623 1165 1626
rect 1154 1566 1157 1623
rect 1154 1563 1165 1566
rect 1114 1533 1141 1536
rect 1106 1443 1109 1516
rect 1114 1506 1117 1533
rect 1114 1503 1125 1506
rect 1130 1503 1133 1526
rect 1146 1503 1149 1516
rect 1106 1413 1109 1436
rect 986 1356 989 1376
rect 986 1353 993 1356
rect 962 1206 965 1326
rect 990 1306 993 1353
rect 1002 1313 1005 1336
rect 1034 1326 1037 1346
rect 1026 1323 1037 1326
rect 986 1303 993 1306
rect 962 1203 969 1206
rect 946 1123 949 1136
rect 954 1106 957 1196
rect 930 1103 941 1106
rect 938 1026 941 1103
rect 930 1023 941 1026
rect 950 1103 957 1106
rect 950 1026 953 1103
rect 966 1096 969 1203
rect 978 1133 981 1226
rect 986 1193 989 1303
rect 1026 1246 1029 1323
rect 1026 1243 1037 1246
rect 994 1123 997 1206
rect 1010 1203 1013 1226
rect 1034 1213 1037 1243
rect 1042 1213 1045 1386
rect 1050 1293 1053 1336
rect 1066 1313 1069 1396
rect 1082 1316 1085 1386
rect 1090 1323 1093 1376
rect 1074 1313 1085 1316
rect 1082 1293 1085 1306
rect 1058 1203 1061 1226
rect 1098 1213 1101 1316
rect 1122 1223 1125 1503
rect 1130 1413 1141 1416
rect 1130 1393 1133 1406
rect 1146 1393 1149 1446
rect 1154 1413 1157 1546
rect 1162 1406 1165 1563
rect 1154 1403 1165 1406
rect 1154 1216 1157 1403
rect 1170 1396 1173 1626
rect 1178 1583 1181 1640
rect 1202 1563 1205 1640
rect 1218 1533 1221 1626
rect 1226 1553 1229 1640
rect 1242 1563 1245 1640
rect 1258 1613 1261 1640
rect 1202 1506 1205 1526
rect 1202 1503 1213 1506
rect 1162 1393 1173 1396
rect 1178 1373 1181 1436
rect 1186 1366 1189 1436
rect 1210 1416 1213 1503
rect 1178 1363 1189 1366
rect 1202 1413 1213 1416
rect 1226 1413 1229 1546
rect 1274 1543 1277 1640
rect 1242 1503 1245 1526
rect 1162 1303 1165 1326
rect 1178 1323 1181 1363
rect 1146 1213 1157 1216
rect 1178 1213 1181 1236
rect 1018 1146 1021 1186
rect 1010 1143 1021 1146
rect 962 1093 969 1096
rect 1010 1096 1013 1143
rect 1042 1133 1045 1186
rect 1066 1173 1069 1206
rect 1146 1166 1149 1213
rect 1162 1183 1165 1206
rect 1146 1163 1157 1166
rect 1066 1133 1069 1156
rect 1010 1093 1021 1096
rect 950 1023 957 1026
rect 930 1003 933 1023
rect 954 943 957 1023
rect 962 936 965 1093
rect 978 1023 981 1036
rect 1018 1016 1021 1093
rect 1018 1013 1037 1016
rect 978 993 981 1006
rect 898 853 917 856
rect 794 773 801 776
rect 842 773 845 806
rect 914 776 917 853
rect 930 803 933 936
rect 954 933 965 936
rect 986 933 989 946
rect 1034 933 1037 1013
rect 1050 993 1053 1016
rect 1098 993 1101 1106
rect 1114 1013 1117 1126
rect 1114 966 1117 1006
rect 1106 963 1117 966
rect 706 733 717 736
rect 794 723 797 773
rect 850 713 853 736
rect 610 693 621 696
rect 562 603 565 616
rect 578 613 581 626
rect 482 493 501 496
rect 570 456 573 566
rect 554 453 573 456
rect 426 366 429 396
rect 442 383 445 416
rect 466 413 469 426
rect 474 383 477 416
rect 506 413 509 426
rect 410 363 429 366
rect 410 286 413 363
rect 482 333 485 346
rect 514 333 517 346
rect 410 283 421 286
rect 322 103 325 116
rect 330 113 333 126
rect 354 103 357 116
rect 418 13 421 283
rect 434 213 453 216
rect 458 203 461 326
rect 538 276 541 326
rect 530 273 541 276
rect 530 213 533 273
rect 554 223 557 453
rect 586 343 589 576
rect 594 523 597 566
rect 610 563 613 693
rect 618 603 621 626
rect 658 613 661 626
rect 810 623 829 626
rect 634 563 637 606
rect 714 593 717 616
rect 722 603 725 616
rect 810 613 813 623
rect 826 613 829 623
rect 682 533 685 576
rect 666 513 669 526
rect 602 316 605 346
rect 618 333 621 416
rect 698 413 701 436
rect 634 323 637 366
rect 602 313 613 316
rect 586 276 589 296
rect 578 273 589 276
rect 530 193 533 206
rect 482 123 485 136
rect 554 133 557 216
rect 578 196 581 273
rect 610 266 613 313
rect 658 306 661 326
rect 602 263 613 266
rect 650 303 661 306
rect 602 203 605 263
rect 650 236 653 303
rect 666 246 669 396
rect 706 346 709 416
rect 714 356 717 526
rect 722 393 725 406
rect 730 393 733 406
rect 714 353 725 356
rect 706 343 717 346
rect 666 243 673 246
rect 650 233 661 236
rect 626 203 629 216
rect 658 213 661 233
rect 578 193 589 196
rect 634 193 637 206
rect 586 133 589 193
rect 658 133 661 196
rect 670 146 673 243
rect 682 223 685 236
rect 690 223 693 326
rect 698 323 701 336
rect 714 333 717 343
rect 722 333 725 353
rect 722 313 725 326
rect 738 296 741 416
rect 746 366 749 606
rect 754 526 757 606
rect 810 593 813 606
rect 834 593 837 616
rect 842 603 845 616
rect 850 613 853 706
rect 866 603 869 776
rect 906 773 917 776
rect 890 713 893 726
rect 906 666 909 773
rect 890 663 909 666
rect 890 623 893 663
rect 946 626 949 806
rect 962 786 965 926
rect 994 923 1005 926
rect 1010 913 1013 926
rect 1026 903 1029 926
rect 1042 913 1045 926
rect 1010 813 1013 836
rect 954 733 957 786
rect 962 783 973 786
rect 930 623 949 626
rect 754 523 761 526
rect 758 466 761 523
rect 754 463 761 466
rect 754 393 757 463
rect 770 443 773 526
rect 778 506 781 526
rect 778 503 789 506
rect 786 436 789 503
rect 778 433 789 436
rect 746 363 757 366
rect 730 293 741 296
rect 730 246 733 293
rect 730 243 741 246
rect 666 143 673 146
rect 546 113 549 126
rect 554 93 557 116
rect 450 0 453 16
rect 562 0 565 126
rect 570 113 573 126
rect 626 103 629 116
rect 634 103 637 126
rect 642 93 645 126
rect 650 113 653 126
rect 658 103 661 116
rect 642 0 645 86
rect 666 83 669 143
rect 674 93 677 126
rect 682 123 685 136
rect 698 133 701 236
rect 706 213 709 236
rect 738 133 741 243
rect 754 166 757 363
rect 778 216 781 433
rect 794 393 797 416
rect 818 403 821 416
rect 834 413 837 526
rect 850 403 853 416
rect 858 413 861 536
rect 874 513 877 606
rect 898 523 909 526
rect 818 326 821 336
rect 794 323 821 326
rect 778 213 785 216
rect 746 163 757 166
rect 746 143 749 163
rect 738 106 741 126
rect 746 116 749 136
rect 746 113 757 116
rect 730 103 741 106
rect 730 16 733 103
rect 730 13 741 16
rect 738 0 741 13
rect 754 0 757 113
rect 770 0 773 146
rect 782 126 785 213
rect 782 123 789 126
rect 794 123 797 323
rect 810 293 813 306
rect 818 286 821 316
rect 810 283 821 286
rect 810 146 813 283
rect 818 203 821 236
rect 826 213 829 226
rect 810 143 821 146
rect 802 123 805 136
rect 818 123 821 143
rect 874 123 885 126
rect 786 106 789 123
rect 786 103 797 106
rect 794 16 797 103
rect 890 93 893 406
rect 898 396 901 406
rect 906 403 909 436
rect 914 413 917 426
rect 922 396 925 416
rect 930 403 933 623
rect 954 613 957 636
rect 970 613 973 783
rect 986 776 989 806
rect 982 773 989 776
rect 982 726 985 773
rect 994 733 997 806
rect 1026 796 1029 826
rect 1042 806 1045 896
rect 1066 893 1069 936
rect 1090 853 1093 926
rect 1098 923 1101 936
rect 1106 856 1109 963
rect 1106 853 1113 856
rect 1066 813 1069 846
rect 1090 823 1093 836
rect 1042 803 1053 806
rect 1026 793 1037 796
rect 982 723 989 726
rect 986 636 989 723
rect 986 633 997 636
rect 938 533 941 606
rect 954 593 957 606
rect 978 593 981 626
rect 994 586 997 633
rect 1010 613 1013 736
rect 1018 693 1021 726
rect 1034 723 1037 793
rect 1050 756 1053 803
rect 1046 753 1053 756
rect 986 583 997 586
rect 946 523 949 546
rect 954 436 957 526
rect 986 456 989 583
rect 1010 513 1013 606
rect 1026 603 1029 616
rect 1034 536 1037 716
rect 1046 636 1049 753
rect 1058 713 1061 736
rect 1082 733 1085 806
rect 1110 776 1113 853
rect 1106 773 1113 776
rect 1082 703 1085 726
rect 1106 723 1109 773
rect 1122 706 1125 996
rect 1146 946 1149 1146
rect 1154 1123 1157 1163
rect 1170 1143 1173 1206
rect 1186 1136 1189 1336
rect 1202 1333 1205 1413
rect 1210 1373 1213 1406
rect 1194 1303 1197 1326
rect 1194 1213 1197 1226
rect 1170 1133 1189 1136
rect 1154 1013 1157 1026
rect 1170 1013 1173 1133
rect 1178 1123 1197 1126
rect 1178 1106 1181 1123
rect 1178 1103 1189 1106
rect 1186 1046 1189 1103
rect 1178 1043 1189 1046
rect 1178 1023 1181 1043
rect 1202 1023 1205 1116
rect 1170 953 1173 1006
rect 1178 1003 1181 1016
rect 1146 943 1157 946
rect 1154 896 1157 943
rect 1146 893 1157 896
rect 1146 836 1149 893
rect 1138 833 1149 836
rect 1138 816 1141 833
rect 1134 813 1141 816
rect 1134 746 1137 813
rect 1134 743 1141 746
rect 1114 703 1125 706
rect 1042 633 1049 636
rect 1042 596 1045 633
rect 1050 603 1053 616
rect 1042 593 1053 596
rect 1050 543 1053 593
rect 1114 543 1117 703
rect 1026 533 1037 536
rect 986 453 997 456
rect 946 433 957 436
rect 978 433 981 446
rect 898 393 925 396
rect 914 193 917 356
rect 922 343 925 393
rect 922 323 925 336
rect 930 333 933 396
rect 938 323 941 426
rect 946 353 949 433
rect 954 346 957 416
rect 978 406 981 426
rect 962 403 981 406
rect 962 363 965 403
rect 994 396 997 453
rect 1010 413 1013 426
rect 1018 396 1021 436
rect 1026 423 1029 533
rect 1034 506 1037 526
rect 1122 523 1125 626
rect 1130 516 1133 726
rect 1138 613 1141 743
rect 1146 546 1149 826
rect 1162 733 1165 826
rect 1170 803 1173 926
rect 1194 913 1197 1016
rect 1218 1013 1221 1326
rect 1242 1293 1245 1326
rect 1242 1223 1245 1246
rect 1250 1203 1253 1376
rect 1258 1323 1261 1426
rect 1266 1373 1269 1406
rect 1282 1393 1285 1566
rect 1290 1533 1293 1640
rect 1306 1623 1309 1640
rect 1298 1596 1301 1616
rect 1298 1593 1305 1596
rect 1302 1526 1305 1593
rect 1298 1523 1305 1526
rect 1314 1523 1317 1606
rect 1338 1566 1341 1586
rect 1330 1563 1341 1566
rect 1298 1456 1301 1523
rect 1330 1486 1333 1563
rect 1354 1526 1357 1640
rect 1362 1533 1365 1546
rect 1354 1523 1365 1526
rect 1354 1503 1357 1516
rect 1330 1483 1341 1486
rect 1294 1453 1301 1456
rect 1294 1386 1297 1453
rect 1314 1413 1317 1426
rect 1338 1413 1341 1483
rect 1362 1456 1365 1523
rect 1378 1503 1381 1526
rect 1386 1496 1389 1546
rect 1434 1533 1437 1556
rect 1450 1533 1453 1640
rect 1474 1566 1477 1640
rect 1470 1563 1477 1566
rect 1354 1453 1365 1456
rect 1378 1493 1389 1496
rect 1294 1383 1301 1386
rect 1266 1296 1269 1366
rect 1298 1363 1301 1383
rect 1322 1376 1325 1406
rect 1314 1373 1325 1376
rect 1354 1376 1357 1453
rect 1370 1423 1373 1436
rect 1354 1373 1365 1376
rect 1378 1373 1381 1493
rect 1394 1413 1397 1436
rect 1410 1416 1413 1526
rect 1402 1413 1413 1416
rect 1418 1413 1429 1416
rect 1442 1413 1445 1436
rect 1402 1406 1405 1413
rect 1394 1403 1405 1406
rect 1314 1333 1317 1373
rect 1274 1313 1277 1326
rect 1306 1303 1309 1316
rect 1330 1303 1333 1326
rect 1362 1306 1365 1373
rect 1362 1303 1373 1306
rect 1266 1293 1277 1296
rect 1274 1236 1277 1293
rect 1266 1233 1277 1236
rect 1266 1183 1269 1233
rect 1314 1223 1317 1236
rect 1322 1203 1325 1216
rect 1338 1213 1341 1246
rect 1266 1133 1269 1156
rect 1346 1146 1349 1256
rect 1354 1213 1357 1296
rect 1370 1256 1373 1303
rect 1394 1276 1397 1403
rect 1418 1393 1421 1406
rect 1450 1383 1453 1406
rect 1458 1393 1461 1526
rect 1470 1486 1473 1563
rect 1546 1556 1549 1640
rect 1546 1553 1557 1556
rect 1470 1483 1477 1486
rect 1402 1333 1405 1346
rect 1418 1336 1421 1366
rect 1410 1333 1421 1336
rect 1410 1306 1413 1326
rect 1362 1253 1373 1256
rect 1386 1273 1397 1276
rect 1406 1303 1413 1306
rect 1338 1143 1349 1146
rect 1234 1056 1237 1126
rect 1250 1103 1253 1116
rect 1314 1113 1317 1126
rect 1230 1053 1237 1056
rect 1202 923 1205 956
rect 1210 936 1213 1006
rect 1230 966 1233 1053
rect 1338 1016 1341 1143
rect 1362 1136 1365 1253
rect 1370 1213 1373 1236
rect 1386 1213 1389 1273
rect 1354 1133 1365 1136
rect 1354 1096 1357 1116
rect 1350 1093 1357 1096
rect 1350 1036 1353 1093
rect 1350 1033 1357 1036
rect 1250 976 1253 1016
rect 1298 983 1301 1006
rect 1242 973 1253 976
rect 1230 963 1237 966
rect 1234 943 1237 963
rect 1210 933 1221 936
rect 1242 933 1245 973
rect 1250 926 1253 946
rect 1258 933 1261 956
rect 1178 813 1189 816
rect 1210 813 1213 926
rect 1218 923 1237 926
rect 1242 923 1253 926
rect 1218 896 1221 916
rect 1242 913 1245 923
rect 1218 893 1237 896
rect 1178 733 1181 746
rect 1154 646 1157 726
rect 1170 666 1173 726
rect 1186 723 1189 813
rect 1202 723 1205 736
rect 1210 723 1213 806
rect 1234 756 1237 893
rect 1218 753 1237 756
rect 1170 663 1181 666
rect 1154 643 1165 646
rect 1162 576 1165 643
rect 1178 613 1181 663
rect 1194 613 1197 626
rect 1218 613 1221 753
rect 1250 613 1253 736
rect 1266 733 1269 976
rect 1306 933 1309 976
rect 1314 926 1317 1016
rect 1338 1013 1349 1016
rect 1322 993 1325 1006
rect 1346 993 1349 1013
rect 1354 1003 1357 1033
rect 1362 1023 1365 1126
rect 1370 1103 1373 1116
rect 1306 923 1317 926
rect 1274 823 1277 846
rect 1306 746 1309 923
rect 1314 903 1317 916
rect 1298 743 1309 746
rect 1274 703 1277 716
rect 1186 593 1189 606
rect 1282 593 1285 616
rect 1298 596 1301 743
rect 1306 723 1309 736
rect 1322 733 1325 796
rect 1330 783 1333 816
rect 1346 813 1349 946
rect 1362 933 1365 976
rect 1378 966 1381 1156
rect 1394 1113 1397 1226
rect 1406 1216 1409 1303
rect 1418 1253 1421 1333
rect 1434 1313 1437 1336
rect 1442 1333 1445 1346
rect 1474 1333 1477 1483
rect 1490 1346 1493 1426
rect 1498 1403 1501 1526
rect 1538 1523 1541 1536
rect 1482 1343 1493 1346
rect 1514 1346 1517 1416
rect 1522 1363 1525 1406
rect 1530 1383 1533 1416
rect 1554 1413 1557 1553
rect 1562 1523 1565 1640
rect 1634 1453 1637 1526
rect 1658 1446 1661 1536
rect 1698 1533 1701 1556
rect 1682 1496 1685 1516
rect 1642 1443 1661 1446
rect 1674 1493 1685 1496
rect 1618 1403 1621 1416
rect 1514 1343 1533 1346
rect 1482 1316 1485 1343
rect 1490 1333 1509 1336
rect 1506 1323 1509 1333
rect 1482 1313 1509 1316
rect 1506 1223 1509 1313
rect 1530 1236 1533 1343
rect 1562 1313 1565 1326
rect 1610 1286 1613 1346
rect 1626 1333 1629 1386
rect 1642 1343 1645 1443
rect 1674 1436 1677 1493
rect 1674 1433 1685 1436
rect 1658 1333 1661 1406
rect 1666 1363 1669 1406
rect 1610 1283 1629 1286
rect 1514 1233 1533 1236
rect 1402 1213 1409 1216
rect 1402 1123 1405 1213
rect 1410 1183 1413 1206
rect 1426 1153 1429 1206
rect 1474 1163 1477 1216
rect 1506 1206 1509 1216
rect 1514 1213 1517 1233
rect 1506 1203 1517 1206
rect 1442 1056 1445 1146
rect 1442 1053 1449 1056
rect 1426 993 1429 1016
rect 1446 1006 1449 1053
rect 1458 1013 1461 1136
rect 1466 1106 1469 1136
rect 1506 1133 1509 1166
rect 1514 1133 1517 1203
rect 1522 1133 1525 1216
rect 1530 1183 1533 1216
rect 1602 1213 1605 1236
rect 1474 1123 1485 1126
rect 1466 1103 1473 1106
rect 1470 1036 1473 1103
rect 1466 1033 1473 1036
rect 1466 1006 1469 1033
rect 1442 1003 1449 1006
rect 1458 1003 1469 1006
rect 1394 966 1397 986
rect 1442 983 1445 1003
rect 1378 963 1389 966
rect 1394 963 1401 966
rect 1370 913 1373 926
rect 1386 876 1389 963
rect 1382 873 1389 876
rect 1354 823 1357 856
rect 1346 793 1349 806
rect 1370 733 1373 816
rect 1382 746 1385 873
rect 1398 866 1401 963
rect 1410 933 1413 946
rect 1458 933 1461 1003
rect 1474 996 1477 1016
rect 1482 1003 1485 1123
rect 1498 1096 1501 1126
rect 1514 1113 1517 1126
rect 1498 1093 1509 1096
rect 1506 1026 1509 1093
rect 1562 1056 1565 1076
rect 1554 1053 1565 1056
rect 1506 1023 1525 1026
rect 1466 993 1477 996
rect 1410 903 1413 926
rect 1466 916 1469 993
rect 1462 913 1469 916
rect 1394 863 1401 866
rect 1394 763 1397 863
rect 1462 846 1465 913
rect 1462 843 1469 846
rect 1382 743 1389 746
rect 1330 693 1333 716
rect 1370 706 1373 726
rect 1362 703 1373 706
rect 1330 603 1333 636
rect 1298 593 1317 596
rect 1162 573 1173 576
rect 1146 543 1157 546
rect 1122 513 1133 516
rect 1034 503 1045 506
rect 1042 436 1045 503
rect 1098 436 1101 446
rect 1034 433 1045 436
rect 1090 433 1101 436
rect 986 393 997 396
rect 1010 393 1021 396
rect 1034 396 1037 433
rect 1066 396 1069 416
rect 1034 393 1045 396
rect 946 306 949 346
rect 954 343 961 346
rect 938 303 949 306
rect 938 236 941 303
rect 958 296 961 343
rect 986 306 989 393
rect 1010 336 1013 393
rect 1010 333 1021 336
rect 986 303 997 306
rect 954 293 961 296
rect 938 233 949 236
rect 922 213 925 226
rect 930 123 933 206
rect 946 203 949 233
rect 954 213 957 293
rect 954 193 957 206
rect 954 133 957 146
rect 786 13 797 16
rect 786 0 789 13
rect 874 0 877 26
rect 922 0 925 16
rect 938 0 941 96
rect 970 13 973 296
rect 994 46 997 303
rect 1018 253 1021 333
rect 1026 323 1029 366
rect 1042 326 1045 393
rect 1058 393 1069 396
rect 1058 336 1061 393
rect 1058 333 1069 336
rect 1034 323 1045 326
rect 1018 123 1021 246
rect 1034 213 1037 323
rect 1066 313 1069 333
rect 1074 313 1077 426
rect 1090 403 1093 433
rect 1098 396 1101 426
rect 1122 413 1125 426
rect 1090 393 1101 396
rect 1050 223 1053 306
rect 1058 233 1061 256
rect 1026 153 1029 206
rect 1042 203 1045 216
rect 1082 213 1085 326
rect 1090 303 1093 393
rect 1130 316 1133 513
rect 1138 406 1141 536
rect 1154 466 1157 543
rect 1146 463 1157 466
rect 1146 413 1149 463
rect 1170 446 1173 573
rect 1218 476 1221 546
rect 1266 486 1269 526
rect 1266 483 1277 486
rect 1218 473 1229 476
rect 1154 443 1173 446
rect 1154 413 1157 443
rect 1162 413 1165 426
rect 1226 416 1229 473
rect 1218 413 1229 416
rect 1250 413 1253 436
rect 1266 413 1269 426
rect 1138 403 1149 406
rect 1218 356 1221 413
rect 1218 353 1229 356
rect 1130 313 1141 316
rect 1130 223 1133 246
rect 1034 133 1037 146
rect 1058 123 1061 156
rect 1122 133 1125 206
rect 1146 146 1149 336
rect 1178 313 1181 326
rect 1186 213 1189 336
rect 1202 313 1205 326
rect 1210 323 1213 336
rect 1146 143 1165 146
rect 1162 126 1165 143
rect 1114 113 1117 126
rect 1154 123 1165 126
rect 986 43 997 46
rect 986 23 989 43
rect 1154 0 1157 123
rect 1194 116 1197 136
rect 1202 123 1205 206
rect 1210 116 1213 126
rect 1226 123 1229 353
rect 1242 333 1245 406
rect 1250 243 1253 406
rect 1274 403 1277 483
rect 1282 413 1285 436
rect 1314 403 1317 593
rect 1362 556 1365 703
rect 1378 603 1381 726
rect 1386 716 1389 743
rect 1410 733 1413 806
rect 1466 803 1469 843
rect 1474 823 1477 936
rect 1482 813 1485 926
rect 1490 766 1493 946
rect 1498 923 1501 976
rect 1506 933 1509 1016
rect 1514 993 1517 1006
rect 1522 983 1525 1023
rect 1530 973 1533 1006
rect 1554 986 1557 1053
rect 1578 1036 1581 1156
rect 1626 1153 1629 1283
rect 1658 1226 1661 1326
rect 1674 1246 1677 1416
rect 1682 1323 1685 1433
rect 1690 1423 1693 1526
rect 1698 1403 1701 1456
rect 1674 1243 1685 1246
rect 1658 1223 1669 1226
rect 1642 1183 1645 1206
rect 1674 1203 1677 1236
rect 1626 1123 1629 1146
rect 1682 1136 1685 1243
rect 1690 1216 1693 1366
rect 1690 1213 1701 1216
rect 1698 1203 1701 1213
rect 1674 1133 1685 1136
rect 1698 1133 1701 1146
rect 1674 1073 1677 1133
rect 1690 1123 1701 1126
rect 1706 1123 1709 1136
rect 1714 1116 1717 1326
rect 1706 1113 1717 1116
rect 1706 1096 1709 1113
rect 1722 1096 1725 1136
rect 1698 1093 1709 1096
rect 1718 1093 1725 1096
rect 1698 1036 1701 1093
rect 1578 1033 1589 1036
rect 1698 1033 1709 1036
rect 1554 983 1565 986
rect 1506 916 1509 926
rect 1498 913 1509 916
rect 1498 813 1501 913
rect 1506 833 1509 846
rect 1514 836 1517 936
rect 1562 933 1565 983
rect 1586 973 1589 1033
rect 1634 1003 1637 1016
rect 1626 933 1629 996
rect 1634 933 1645 936
rect 1634 926 1637 933
rect 1514 833 1525 836
rect 1506 823 1517 826
rect 1522 806 1525 833
rect 1514 803 1525 806
rect 1530 803 1533 846
rect 1546 813 1549 876
rect 1570 813 1573 926
rect 1594 873 1597 926
rect 1626 923 1637 926
rect 1386 713 1397 716
rect 1394 656 1397 713
rect 1386 653 1397 656
rect 1386 633 1389 653
rect 1362 553 1373 556
rect 1370 533 1373 553
rect 1386 533 1389 616
rect 1402 523 1405 626
rect 1418 523 1421 726
rect 1426 603 1429 626
rect 1434 613 1437 726
rect 1442 713 1445 736
rect 1458 733 1461 766
rect 1490 763 1501 766
rect 1490 733 1493 756
rect 1498 746 1501 763
rect 1498 743 1505 746
rect 1466 723 1485 726
rect 1442 593 1445 606
rect 1330 403 1333 426
rect 1274 333 1285 336
rect 1242 203 1245 216
rect 1282 193 1285 326
rect 1290 323 1293 346
rect 1290 303 1293 316
rect 1298 313 1301 336
rect 1362 223 1365 336
rect 1370 333 1373 346
rect 1362 213 1373 216
rect 1282 123 1285 146
rect 1306 143 1309 206
rect 1370 143 1373 156
rect 1194 113 1213 116
rect 1194 0 1197 113
rect 1306 103 1309 136
rect 1378 133 1381 236
rect 1394 206 1397 516
rect 1434 513 1437 536
rect 1450 523 1453 616
rect 1458 503 1461 716
rect 1466 703 1469 716
rect 1466 613 1469 626
rect 1466 533 1469 596
rect 1474 526 1477 606
rect 1490 546 1493 726
rect 1502 636 1505 743
rect 1514 723 1517 803
rect 1522 763 1525 796
rect 1502 633 1509 636
rect 1506 616 1509 633
rect 1514 623 1517 706
rect 1506 613 1517 616
rect 1514 603 1517 613
rect 1522 593 1525 736
rect 1538 713 1541 806
rect 1562 733 1565 786
rect 1594 763 1597 816
rect 1602 796 1605 836
rect 1626 813 1629 923
rect 1634 813 1637 826
rect 1642 796 1645 846
rect 1650 813 1653 926
rect 1658 833 1661 986
rect 1666 933 1669 1006
rect 1674 993 1677 1006
rect 1674 923 1677 936
rect 1682 933 1685 1016
rect 1674 823 1677 846
rect 1602 793 1613 796
rect 1578 733 1581 756
rect 1554 603 1557 726
rect 1570 693 1573 726
rect 1594 693 1597 716
rect 1610 686 1613 793
rect 1634 793 1645 796
rect 1650 793 1653 806
rect 1634 703 1637 793
rect 1658 746 1661 816
rect 1666 813 1677 816
rect 1690 803 1693 976
rect 1698 923 1701 1016
rect 1706 1013 1709 1033
rect 1718 1026 1721 1093
rect 1714 1023 1721 1026
rect 1714 996 1717 1023
rect 1710 993 1717 996
rect 1710 856 1713 993
rect 1710 853 1717 856
rect 1714 776 1717 853
rect 1722 806 1725 1016
rect 1730 1013 1733 1216
rect 1738 1116 1741 1136
rect 1738 1113 1749 1116
rect 1746 1036 1749 1113
rect 1738 1033 1749 1036
rect 1730 966 1733 1006
rect 1738 983 1741 1033
rect 1730 963 1741 966
rect 1738 866 1741 963
rect 1754 923 1757 1006
rect 1730 863 1741 866
rect 1730 813 1733 863
rect 1770 813 1773 826
rect 1722 803 1733 806
rect 1698 773 1717 776
rect 1658 743 1669 746
rect 1658 726 1661 736
rect 1642 723 1661 726
rect 1666 723 1669 743
rect 1698 733 1701 773
rect 1698 723 1717 726
rect 1602 683 1613 686
rect 1594 576 1597 596
rect 1590 573 1597 576
rect 1490 543 1501 546
rect 1466 523 1477 526
rect 1426 403 1445 406
rect 1434 333 1437 356
rect 1442 323 1445 403
rect 1450 353 1453 406
rect 1458 346 1461 406
rect 1450 343 1461 346
rect 1450 316 1453 343
rect 1466 326 1469 523
rect 1490 516 1493 536
rect 1486 513 1493 516
rect 1442 313 1453 316
rect 1462 323 1469 326
rect 1442 266 1445 313
rect 1442 263 1453 266
rect 1394 203 1405 206
rect 1386 133 1389 156
rect 1402 146 1405 203
rect 1450 196 1453 263
rect 1462 256 1465 323
rect 1462 253 1469 256
rect 1458 223 1461 236
rect 1466 213 1469 253
rect 1474 206 1477 506
rect 1486 436 1489 513
rect 1486 433 1493 436
rect 1482 393 1485 416
rect 1490 386 1493 433
rect 1498 413 1501 543
rect 1506 516 1509 536
rect 1506 513 1513 516
rect 1510 436 1513 513
rect 1522 496 1525 536
rect 1530 513 1533 526
rect 1554 523 1557 536
rect 1578 506 1581 536
rect 1570 503 1581 506
rect 1522 493 1533 496
rect 1530 436 1533 493
rect 1506 433 1513 436
rect 1522 433 1533 436
rect 1506 386 1509 433
rect 1522 413 1525 433
rect 1482 383 1493 386
rect 1498 383 1509 386
rect 1522 403 1533 406
rect 1482 316 1485 383
rect 1490 333 1493 356
rect 1498 323 1501 383
rect 1482 313 1489 316
rect 1486 246 1489 313
rect 1394 143 1405 146
rect 1442 193 1453 196
rect 1458 203 1477 206
rect 1482 243 1489 246
rect 1394 123 1397 143
rect 1434 116 1437 136
rect 1442 123 1445 193
rect 1450 133 1453 146
rect 1458 123 1461 203
rect 1482 143 1485 243
rect 1466 123 1469 136
rect 1490 123 1493 226
rect 1506 213 1509 336
rect 1522 333 1525 403
rect 1570 366 1573 503
rect 1590 486 1593 573
rect 1602 533 1605 683
rect 1626 593 1629 616
rect 1642 546 1645 616
rect 1658 613 1661 716
rect 1682 653 1685 716
rect 1690 703 1693 716
rect 1722 606 1725 796
rect 1730 733 1733 803
rect 1730 723 1749 726
rect 1730 703 1733 716
rect 1618 533 1621 546
rect 1626 543 1645 546
rect 1626 523 1629 543
rect 1602 496 1605 516
rect 1634 513 1637 526
rect 1642 496 1645 536
rect 1602 493 1613 496
rect 1590 483 1597 486
rect 1570 363 1581 366
rect 1522 236 1525 326
rect 1538 316 1541 336
rect 1570 323 1573 346
rect 1578 333 1581 363
rect 1586 323 1589 356
rect 1594 333 1597 483
rect 1610 436 1613 493
rect 1602 433 1613 436
rect 1634 493 1645 496
rect 1634 436 1637 493
rect 1650 446 1653 606
rect 1682 593 1685 606
rect 1722 603 1733 606
rect 1666 516 1669 536
rect 1722 533 1725 596
rect 1666 513 1677 516
rect 1698 513 1701 526
rect 1674 446 1677 513
rect 1650 443 1657 446
rect 1634 433 1645 436
rect 1602 403 1605 433
rect 1610 403 1613 416
rect 1642 413 1645 433
rect 1618 393 1621 406
rect 1634 326 1637 406
rect 1642 393 1645 406
rect 1654 396 1657 443
rect 1666 443 1677 446
rect 1666 406 1669 443
rect 1674 413 1677 426
rect 1714 423 1717 516
rect 1722 496 1725 526
rect 1730 523 1733 603
rect 1746 556 1749 626
rect 1754 613 1757 726
rect 1738 553 1749 556
rect 1738 516 1741 553
rect 1730 513 1741 516
rect 1722 493 1733 496
rect 1730 436 1733 493
rect 1754 473 1757 546
rect 1722 433 1733 436
rect 1722 413 1725 433
rect 1770 413 1773 476
rect 1666 403 1677 406
rect 1654 393 1669 396
rect 1634 323 1653 326
rect 1538 313 1549 316
rect 1546 246 1549 313
rect 1650 306 1653 323
rect 1514 233 1525 236
rect 1538 243 1549 246
rect 1642 303 1653 306
rect 1658 306 1661 336
rect 1666 323 1669 393
rect 1674 333 1677 403
rect 1658 303 1669 306
rect 1642 246 1645 303
rect 1666 246 1669 303
rect 1642 243 1653 246
rect 1514 206 1517 233
rect 1530 213 1533 226
rect 1506 203 1517 206
rect 1538 203 1541 243
rect 1506 133 1509 203
rect 1546 193 1549 226
rect 1586 203 1589 236
rect 1650 226 1653 243
rect 1634 213 1637 226
rect 1642 223 1653 226
rect 1658 243 1669 246
rect 1658 223 1661 243
rect 1642 213 1645 223
rect 1618 203 1637 206
rect 1530 133 1533 146
rect 1434 113 1453 116
rect 1530 113 1533 126
rect 1538 113 1541 126
rect 1570 123 1573 146
rect 1450 0 1453 113
rect 1618 103 1621 146
rect 1634 133 1637 203
rect 1642 193 1645 206
rect 1650 203 1653 216
rect 1658 133 1661 206
rect 1666 133 1669 216
rect 1674 203 1677 216
rect 1690 133 1693 406
rect 1770 366 1773 386
rect 1762 363 1773 366
rect 1762 266 1765 363
rect 1762 263 1773 266
rect 1714 213 1717 226
rect 1714 123 1717 136
rect 1770 123 1773 263
rect 1778 213 1781 436
rect 1791 37 1811 1603
rect 1815 13 1835 1627
<< metal3 >>
rect 753 1622 870 1627
rect 889 1622 966 1627
rect 1089 1622 1174 1627
rect 1217 1622 1310 1627
rect 1257 1612 1302 1617
rect 1089 1602 1126 1607
rect 1177 1602 1318 1607
rect 1009 1582 1182 1587
rect 1201 1582 1342 1587
rect 729 1572 822 1577
rect 513 1562 614 1567
rect 817 1562 854 1567
rect 1065 1562 1206 1567
rect 1241 1562 1286 1567
rect 385 1552 454 1557
rect 385 1547 390 1552
rect 161 1542 390 1547
rect 449 1547 454 1552
rect 513 1547 518 1562
rect 609 1557 614 1562
rect 609 1552 638 1557
rect 1201 1552 1230 1557
rect 1433 1552 1702 1557
rect 449 1542 518 1547
rect 529 1542 750 1547
rect 841 1542 942 1547
rect 953 1542 974 1547
rect 1105 1542 1158 1547
rect 401 1532 438 1537
rect 545 1532 574 1537
rect 1049 1522 1134 1527
rect 1201 1522 1206 1552
rect 1225 1542 1278 1547
rect 1361 1542 1390 1547
rect 1537 1522 1662 1527
rect 137 1512 190 1517
rect 273 1512 302 1517
rect 441 1512 542 1517
rect 801 1512 854 1517
rect 937 1512 1022 1517
rect 489 1502 590 1507
rect 1145 1502 1246 1507
rect 1353 1502 1382 1507
rect 81 1492 166 1497
rect 689 1452 838 1457
rect 1633 1452 1702 1457
rect 729 1442 758 1447
rect 753 1437 758 1442
rect 817 1442 1054 1447
rect 1105 1442 1150 1447
rect 817 1437 822 1442
rect 753 1432 822 1437
rect 841 1432 878 1437
rect 1105 1432 1182 1437
rect 1369 1432 1398 1437
rect 1409 1432 1446 1437
rect 105 1422 270 1427
rect 601 1422 710 1427
rect 337 1412 414 1417
rect 745 1412 854 1417
rect 985 1412 1046 1417
rect 337 1407 342 1412
rect 225 1402 342 1407
rect 409 1407 414 1412
rect 409 1402 598 1407
rect 617 1402 646 1407
rect 593 1397 598 1402
rect 641 1397 646 1402
rect 769 1402 806 1407
rect 769 1397 774 1402
rect 593 1392 614 1397
rect 641 1392 774 1397
rect 833 1392 1022 1397
rect 161 1382 454 1387
rect 793 1382 966 1387
rect 1041 1382 1046 1412
rect 1089 1397 1094 1417
rect 1065 1392 1094 1397
rect 1105 1412 1142 1417
rect 1313 1412 1422 1417
rect 1105 1387 1110 1412
rect 1161 1402 1262 1407
rect 1617 1402 1662 1407
rect 1161 1397 1166 1402
rect 1129 1392 1166 1397
rect 1257 1397 1262 1402
rect 1257 1392 1286 1397
rect 1417 1392 1462 1397
rect 1081 1382 1110 1387
rect 1449 1382 1630 1387
rect 953 1372 990 1377
rect 1089 1372 1182 1377
rect 1209 1372 1382 1377
rect 153 1362 206 1367
rect 281 1362 406 1367
rect 569 1362 814 1367
rect 929 1362 966 1367
rect 1265 1362 1302 1367
rect 1417 1362 1694 1367
rect 833 1352 854 1357
rect 905 1352 950 1357
rect 137 1342 350 1347
rect 601 1342 822 1347
rect 857 1342 934 1347
rect 545 1332 638 1337
rect 769 1332 854 1337
rect 961 1322 966 1362
rect 1401 1342 1446 1347
rect 1609 1342 1646 1347
rect 1145 1322 1254 1327
rect 1657 1322 1686 1327
rect 1145 1317 1150 1322
rect 169 1312 246 1317
rect 641 1312 750 1317
rect 1001 1312 1150 1317
rect 1249 1317 1254 1322
rect 1249 1312 1278 1317
rect 1433 1312 1566 1317
rect 473 1302 782 1307
rect 1161 1302 1246 1307
rect 1305 1302 1334 1307
rect 177 1292 222 1297
rect 849 1292 886 1297
rect 1049 1292 1086 1297
rect 1241 1292 1398 1297
rect 1345 1252 1422 1257
rect 553 1242 598 1247
rect 1241 1242 1342 1247
rect 529 1232 614 1237
rect 833 1232 894 1237
rect 1177 1232 1254 1237
rect 1313 1232 1374 1237
rect 1601 1232 1678 1237
rect 249 1222 438 1227
rect 513 1222 638 1227
rect 689 1222 838 1227
rect 833 1217 838 1222
rect 905 1222 1014 1227
rect 1057 1222 1198 1227
rect 1393 1222 1662 1227
rect 905 1217 910 1222
rect 449 1212 478 1217
rect 601 1212 630 1217
rect 833 1212 910 1217
rect 473 1207 606 1212
rect 129 1192 198 1197
rect 313 1192 470 1197
rect 561 1192 638 1197
rect 673 1192 806 1197
rect 953 1192 990 1197
rect 673 1187 678 1192
rect 297 1182 342 1187
rect 409 1182 678 1187
rect 697 1182 726 1187
rect 937 1182 1022 1187
rect 1041 1182 1046 1217
rect 1249 1212 1326 1217
rect 1777 1202 1850 1207
rect 1777 1197 1782 1202
rect 1761 1192 1782 1197
rect 1761 1187 1766 1192
rect 1161 1182 1270 1187
rect 1409 1182 1766 1187
rect 337 1172 422 1177
rect 753 1172 926 1177
rect 921 1167 926 1172
rect 1017 1172 1070 1177
rect 1017 1167 1022 1172
rect 921 1162 1022 1167
rect 1473 1162 1510 1167
rect 281 1152 326 1157
rect 321 1147 326 1152
rect 433 1152 574 1157
rect 769 1152 830 1157
rect 1065 1152 1454 1157
rect 1521 1152 1630 1157
rect 433 1147 438 1152
rect 1449 1147 1526 1152
rect 0 1142 206 1147
rect 321 1142 438 1147
rect 641 1142 710 1147
rect 761 1142 862 1147
rect 1041 1142 1070 1147
rect 1145 1142 1174 1147
rect 1625 1142 1702 1147
rect 209 1132 286 1137
rect 865 1132 894 1137
rect 945 1132 982 1137
rect 1465 1132 1518 1137
rect 1705 1132 1742 1137
rect 601 1122 654 1127
rect 817 1122 878 1127
rect 1697 1122 1726 1127
rect 153 1112 238 1117
rect 305 1112 438 1117
rect 1313 1112 1358 1117
rect 1441 1112 1518 1117
rect 217 1102 294 1107
rect 841 1102 1102 1107
rect 1201 1102 1374 1107
rect 345 1092 374 1097
rect 369 1087 374 1092
rect 449 1092 478 1097
rect 449 1087 454 1092
rect 369 1082 454 1087
rect 1561 1072 1678 1077
rect 185 1062 302 1067
rect 185 1057 190 1062
rect 161 1052 190 1057
rect 297 1057 302 1062
rect 297 1052 326 1057
rect 321 1042 350 1047
rect 185 1032 334 1037
rect 705 1032 838 1037
rect 913 1032 982 1037
rect 521 1022 566 1027
rect 705 1022 734 1027
rect 1153 1022 1206 1027
rect 153 1012 254 1017
rect 1113 1012 1182 1017
rect 1697 1012 1734 1017
rect 1633 1002 1670 1007
rect 153 992 182 997
rect 177 987 182 992
rect 265 992 406 997
rect 729 992 774 997
rect 873 992 966 997
rect 977 992 1054 997
rect 1097 992 1126 997
rect 1209 992 1350 997
rect 1425 992 1518 997
rect 1625 992 1678 997
rect 265 987 270 992
rect 177 982 270 987
rect 617 982 790 987
rect 1121 982 1302 987
rect 1393 982 1446 987
rect 1521 982 1742 987
rect 1265 972 1366 977
rect 1497 972 1534 977
rect 1585 972 1694 977
rect 601 962 630 967
rect 1329 957 1430 962
rect 1169 952 1334 957
rect 1425 952 1534 957
rect 1529 947 1534 952
rect 1617 952 1850 957
rect 1617 947 1622 952
rect 249 942 318 947
rect 529 942 622 947
rect 737 942 894 947
rect 953 942 990 947
rect 1233 942 1254 947
rect 1345 942 1414 947
rect 1489 942 1510 947
rect 1529 942 1622 947
rect 0 932 190 937
rect 385 932 414 937
rect 1097 932 1222 937
rect 1641 932 1678 937
rect 225 922 342 927
rect 1001 922 1086 927
rect 1169 922 1374 927
rect 1649 922 1702 927
rect 1081 917 1174 922
rect 353 912 430 917
rect 625 912 726 917
rect 961 912 1046 917
rect 1193 912 1222 917
rect 769 902 902 907
rect 1025 902 1318 907
rect 1409 902 1518 907
rect 1041 892 1070 897
rect 321 872 454 877
rect 321 867 326 872
rect 65 862 326 867
rect 449 867 454 872
rect 1113 872 1294 877
rect 1545 872 1598 877
rect 449 862 534 867
rect 1113 857 1118 872
rect 1089 852 1118 857
rect 1289 857 1294 872
rect 1289 852 1358 857
rect 337 842 438 847
rect 561 842 774 847
rect 1065 842 1278 847
rect 1505 842 1534 847
rect 1641 842 1678 847
rect 185 832 262 837
rect 1009 832 1094 837
rect 1601 832 1662 837
rect 0 822 70 827
rect 81 822 126 827
rect 321 822 430 827
rect 537 822 622 827
rect 961 822 1030 827
rect 1161 822 1510 827
rect 1633 822 1774 827
rect 1345 812 1374 817
rect 1537 812 1574 817
rect 1625 812 1670 817
rect 833 802 910 807
rect 929 802 998 807
rect 833 797 838 802
rect 137 792 206 797
rect 273 792 526 797
rect 273 787 278 792
rect 0 782 126 787
rect 121 777 126 782
rect 217 782 278 787
rect 521 787 526 792
rect 569 792 654 797
rect 569 787 574 792
rect 521 782 574 787
rect 649 787 654 792
rect 697 792 790 797
rect 809 792 838 797
rect 905 797 910 802
rect 905 792 990 797
rect 1081 792 1350 797
rect 1393 792 1518 797
rect 697 787 702 792
rect 649 782 702 787
rect 785 787 790 792
rect 1393 787 1398 792
rect 785 782 958 787
rect 1329 782 1398 787
rect 1513 787 1518 792
rect 1537 787 1542 812
rect 1649 792 1726 797
rect 1513 782 1566 787
rect 217 777 222 782
rect 121 772 222 777
rect 289 772 446 777
rect 585 772 870 777
rect 401 762 678 767
rect 1393 762 1462 767
rect 1521 762 1598 767
rect 529 752 590 757
rect 1489 752 1582 757
rect 153 742 382 747
rect 489 742 566 747
rect 633 742 694 747
rect 1177 742 1214 747
rect 153 737 158 742
rect 0 732 158 737
rect 377 737 382 742
rect 377 732 710 737
rect 1009 732 1086 737
rect 1305 732 1542 737
rect 169 722 270 727
rect 473 722 798 727
rect 1129 722 1302 727
rect 273 712 374 717
rect 537 712 598 717
rect 593 707 598 712
rect 673 712 702 717
rect 849 712 894 717
rect 1033 712 1062 717
rect 673 707 678 712
rect 1297 707 1302 722
rect 1561 722 1638 727
rect 1561 717 1566 722
rect 1417 712 1446 717
rect 1537 712 1566 717
rect 1633 717 1638 722
rect 1633 712 1662 717
rect 441 702 574 707
rect 593 702 678 707
rect 1081 702 1278 707
rect 1297 702 1734 707
rect 1017 692 1070 697
rect 1065 677 1070 692
rect 1225 692 1334 697
rect 1457 692 1598 697
rect 1225 677 1230 692
rect 1065 672 1230 677
rect 1249 672 1278 677
rect 1273 667 1278 672
rect 1345 672 1850 677
rect 1345 667 1350 672
rect 0 662 126 667
rect 1273 662 1350 667
rect 1521 652 1550 657
rect 1545 647 1550 652
rect 1657 652 1686 657
rect 1657 647 1662 652
rect 289 642 430 647
rect 977 642 1214 647
rect 1545 642 1662 647
rect 977 637 982 642
rect 185 632 262 637
rect 953 632 982 637
rect 1209 637 1214 642
rect 1209 632 1390 637
rect 185 627 190 632
rect 161 622 190 627
rect 257 627 262 632
rect 257 622 350 627
rect 473 622 550 627
rect 617 622 662 627
rect 849 622 934 627
rect 1121 622 1198 627
rect 1425 622 1470 627
rect 849 617 854 622
rect 81 612 198 617
rect 329 612 582 617
rect 825 612 854 617
rect 929 617 934 622
rect 929 612 1142 617
rect 241 602 326 607
rect 417 602 446 607
rect 561 602 726 607
rect 841 602 878 607
rect 1009 602 1054 607
rect 713 592 814 597
rect 833 592 862 597
rect 857 587 862 592
rect 929 592 982 597
rect 1185 592 1286 597
rect 1441 592 1526 597
rect 1593 592 1726 597
rect 929 587 934 592
rect 249 582 486 587
rect 857 582 934 587
rect 249 577 254 582
rect 193 572 254 577
rect 481 577 486 582
rect 481 572 686 577
rect 265 562 470 567
rect 465 557 470 562
rect 545 562 638 567
rect 545 557 550 562
rect 113 552 206 557
rect 465 552 550 557
rect 1641 552 1734 557
rect 1641 547 1646 552
rect 337 542 446 547
rect 945 542 1222 547
rect 1617 542 1646 547
rect 1729 547 1734 552
rect 1729 542 1758 547
rect 0 532 102 537
rect 97 527 102 532
rect 201 532 326 537
rect 473 532 510 537
rect 1553 532 1606 537
rect 1641 532 1734 537
rect 201 527 206 532
rect 321 527 438 532
rect 97 522 206 527
rect 433 522 454 527
rect 465 522 486 527
rect 857 522 902 527
rect 1449 522 1534 527
rect 225 512 342 517
rect 665 512 878 517
rect 1433 512 1502 517
rect 1497 507 1502 512
rect 1577 512 1638 517
rect 1697 512 1734 517
rect 1577 507 1582 512
rect 449 502 494 507
rect 1457 502 1478 507
rect 1497 502 1582 507
rect 0 492 86 497
rect 305 492 358 497
rect 257 482 334 487
rect 321 472 350 477
rect 1753 472 1850 477
rect 793 462 958 467
rect 793 447 798 462
rect 769 442 798 447
rect 953 447 958 462
rect 1001 452 1078 457
rect 1001 447 1006 452
rect 953 442 1006 447
rect 1073 447 1078 452
rect 1073 442 1102 447
rect 1657 442 1734 447
rect 1657 437 1662 442
rect 201 432 366 437
rect 697 432 1022 437
rect 1249 432 1286 437
rect 1593 432 1662 437
rect 1729 437 1734 442
rect 1729 432 1850 437
rect 465 422 510 427
rect 913 422 1126 427
rect 1265 422 1334 427
rect 1673 422 1718 427
rect 0 412 270 417
rect 817 412 862 417
rect 1065 412 1166 417
rect 1481 412 1526 417
rect 177 402 214 407
rect 729 402 854 407
rect 889 402 934 407
rect 1529 402 1614 407
rect 249 392 350 397
rect 417 392 758 397
rect 793 392 822 397
rect 817 387 822 392
rect 905 392 934 397
rect 1617 392 1646 397
rect 905 387 910 392
rect 425 382 478 387
rect 817 382 910 387
rect 1769 382 1850 387
rect 0 372 166 377
rect 633 362 1030 367
rect 913 352 950 357
rect 1433 352 1590 357
rect 481 342 590 347
rect 921 342 950 347
rect 1241 342 1294 347
rect 1569 342 1678 347
rect 601 332 718 337
rect 817 332 926 337
rect 1281 332 1422 337
rect 1417 327 1422 332
rect 1481 332 1526 337
rect 1481 327 1486 332
rect 105 322 254 327
rect 697 322 726 327
rect 1177 322 1214 327
rect 1417 322 1486 327
rect 1137 312 1206 317
rect 1281 312 1302 317
rect 1201 307 1206 312
rect 169 302 198 307
rect 193 297 198 302
rect 265 302 350 307
rect 1201 302 1294 307
rect 265 297 270 302
rect 193 292 270 297
rect 585 292 974 297
rect 1017 252 1062 257
rect 777 242 1022 247
rect 1129 242 1254 247
rect 1385 242 1566 247
rect 777 237 782 242
rect 1385 237 1390 242
rect 257 232 366 237
rect 681 232 782 237
rect 953 232 1054 237
rect 1361 232 1390 237
rect 1561 237 1566 242
rect 1561 232 1590 237
rect 345 222 558 227
rect 809 222 926 227
rect 1033 222 1086 227
rect 1457 222 1534 227
rect 1657 222 1718 227
rect 129 212 238 217
rect 625 212 686 217
rect 681 207 686 212
rect 793 212 830 217
rect 945 212 1046 217
rect 1369 212 1470 217
rect 1481 212 1774 217
rect 793 207 798 212
rect 529 202 606 207
rect 681 202 798 207
rect 817 202 982 207
rect 977 197 982 202
rect 1097 202 1126 207
rect 1201 202 1246 207
rect 1473 202 1654 207
rect 1097 197 1102 202
rect 217 192 270 197
rect 633 192 662 197
rect 913 192 958 197
rect 977 192 1102 197
rect 1281 192 1358 197
rect 1353 187 1358 192
rect 1521 192 1646 197
rect 1521 187 1526 192
rect 1353 182 1526 187
rect 1025 152 1062 157
rect 1369 152 1390 157
rect 745 142 774 147
rect 953 142 1230 147
rect 1281 142 1310 147
rect 1449 142 1486 147
rect 1529 142 1574 147
rect 1617 142 1694 147
rect 1441 132 1470 137
rect 1657 132 1718 137
rect 481 122 638 127
rect 649 122 886 127
rect 1225 122 1310 127
rect 1489 122 1534 127
rect 105 112 334 117
rect 545 112 574 117
rect 969 112 1118 117
rect 1449 112 1542 117
rect 321 102 358 107
rect 625 102 662 107
rect 1305 102 1438 107
rect 1433 97 1438 102
rect 1553 102 1622 107
rect 1553 97 1558 102
rect 553 92 678 97
rect 889 92 942 97
rect 1433 92 1558 97
rect 641 82 670 87
rect 873 22 990 27
rect 417 12 454 17
rect 921 12 974 17
use UART_VIA0  UART_VIA0_0
timestamp 1554483974
transform 1 0 24 0 1 1617
box -10 -10 10 10
use M3_M2  M3_M2_0
timestamp 1554483974
transform 1 0 756 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_1
timestamp 1554483974
transform 1 0 868 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_2
timestamp 1554483974
transform 1 0 892 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_3
timestamp 1554483974
transform 1 0 964 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_4
timestamp 1554483974
transform 1 0 1092 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_5
timestamp 1554483974
transform 1 0 1172 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_6
timestamp 1554483974
transform 1 0 1220 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_7
timestamp 1554483974
transform 1 0 1308 0 1 1625
box -3 -3 3 3
use M3_M2  M3_M2_8
timestamp 1554483974
transform 1 0 1260 0 1 1615
box -3 -3 3 3
use M3_M2  M3_M2_9
timestamp 1554483974
transform 1 0 1300 0 1 1615
box -3 -3 3 3
use UART_VIA0  UART_VIA0_2
timestamp 1554483974
transform 1 0 48 0 1 1593
box -10 -10 10 10
use M3_M2  M3_M2_10
timestamp 1554483974
transform 1 0 1092 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_11
timestamp 1554483974
transform 1 0 1124 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_12
timestamp 1554483974
transform 1 0 1180 0 1 1605
box -3 -3 3 3
use M3_M2  M3_M2_13
timestamp 1554483974
transform 1 0 1316 0 1 1605
box -3 -3 3 3
use UART_VIA0  UART_VIA0_1
timestamp 1554483974
transform 1 0 1825 0 1 1617
box -10 -10 10 10
use M3_M2  M3_M2_14
timestamp 1554483974
transform 1 0 1012 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_15
timestamp 1554483974
transform 1 0 1180 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_16
timestamp 1554483974
transform 1 0 1204 0 1 1585
box -3 -3 3 3
use M3_M2  M3_M2_17
timestamp 1554483974
transform 1 0 1340 0 1 1585
box -3 -3 3 3
use UART_VIA0  UART_VIA0_3
timestamp 1554483974
transform 1 0 1801 0 1 1593
box -10 -10 10 10
use UART_VIA1  UART_VIA1_0
timestamp 1554483974
transform 1 0 48 0 1 1570
box -10 -3 10 3
use M3_M2  M3_M2_31
timestamp 1554483974
transform 1 0 164 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_2
timestamp 1554483974
transform 1 0 164 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_26
timestamp 1554483974
transform 1 0 84 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_27
timestamp 1554483974
transform 1 0 140 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_55
timestamp 1554483974
transform 1 0 140 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_73
timestamp 1554483974
transform 1 0 84 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_74
timestamp 1554483974
transform 1 0 164 0 1 1495
box -3 -3 3 3
use M3_M2  M3_M2_56
timestamp 1554483974
transform 1 0 188 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_32
timestamp 1554483974
transform 1 0 204 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_33
timestamp 1554483974
transform 1 0 228 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_3
timestamp 1554483974
transform 1 0 228 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_28
timestamp 1554483974
transform 1 0 276 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_57
timestamp 1554483974
transform 1 0 276 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_58
timestamp 1554483974
transform 1 0 300 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_29
timestamp 1554483974
transform 1 0 356 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_4
timestamp 1554483974
transform 1 0 372 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_0
timestamp 1554483974
transform 1 0 404 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_46
timestamp 1554483974
transform 1 0 404 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_30
timestamp 1554483974
transform 1 0 396 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_47
timestamp 1554483974
transform 1 0 436 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_5
timestamp 1554483974
transform 1 0 444 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_31
timestamp 1554483974
transform 1 0 444 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_32
timestamp 1554483974
transform 1 0 452 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_59
timestamp 1554483974
transform 1 0 444 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_50
timestamp 1554483974
transform 1 0 492 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_66
timestamp 1554483974
transform 1 0 492 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_60
timestamp 1554483974
transform 1 0 516 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_34
timestamp 1554483974
transform 1 0 532 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_6
timestamp 1554483974
transform 1 0 532 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_7
timestamp 1554483974
transform 1 0 540 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_48
timestamp 1554483974
transform 1 0 548 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_33
timestamp 1554483974
transform 1 0 548 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_61
timestamp 1554483974
transform 1 0 540 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_49
timestamp 1554483974
transform 1 0 572 0 1 1535
box -3 -3 3 3
use M2_M1  M2_M1_51
timestamp 1554483974
transform 1 0 564 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_67
timestamp 1554483974
transform 1 0 564 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_68
timestamp 1554483974
transform 1 0 588 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_8
timestamp 1554483974
transform 1 0 604 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_26
timestamp 1554483974
transform 1 0 636 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_9
timestamp 1554483974
transform 1 0 636 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_34
timestamp 1554483974
transform 1 0 684 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_18
timestamp 1554483974
transform 1 0 732 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_35
timestamp 1554483974
transform 1 0 748 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_10
timestamp 1554483974
transform 1 0 748 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_35
timestamp 1554483974
transform 1 0 748 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_19
timestamp 1554483974
transform 1 0 820 0 1 1575
box -3 -3 3 3
use M3_M2  M3_M2_20
timestamp 1554483974
transform 1 0 820 0 1 1565
box -3 -3 3 3
use M2_M1  M2_M1_11
timestamp 1554483974
transform 1 0 804 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_62
timestamp 1554483974
transform 1 0 804 0 1 1515
box -3 -3 3 3
use M3_M2  M3_M2_21
timestamp 1554483974
transform 1 0 852 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_36
timestamp 1554483974
transform 1 0 844 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_12
timestamp 1554483974
transform 1 0 844 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_36
timestamp 1554483974
transform 1 0 836 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_37
timestamp 1554483974
transform 1 0 852 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_63
timestamp 1554483974
transform 1 0 852 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_13
timestamp 1554483974
transform 1 0 900 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_37
timestamp 1554483974
transform 1 0 940 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_38
timestamp 1554483974
transform 1 0 956 0 1 1545
box -3 -3 3 3
use M3_M2  M3_M2_39
timestamp 1554483974
transform 1 0 972 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_14
timestamp 1554483974
transform 1 0 988 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_38
timestamp 1554483974
transform 1 0 908 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_39
timestamp 1554483974
transform 1 0 940 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_64
timestamp 1554483974
transform 1 0 940 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_1
timestamp 1554483974
transform 1 0 1028 0 1 1545
box -2 -2 2 2
use M3_M2  M3_M2_65
timestamp 1554483974
transform 1 0 1020 0 1 1515
box -3 -3 3 3
use M2_M1  M2_M1_15
timestamp 1554483974
transform 1 0 1052 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_40
timestamp 1554483974
transform 1 0 1044 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_50
timestamp 1554483974
transform 1 0 1052 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_22
timestamp 1554483974
transform 1 0 1068 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_40
timestamp 1554483974
transform 1 0 1108 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_52
timestamp 1554483974
transform 1 0 1108 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_51
timestamp 1554483974
transform 1 0 1132 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_41
timestamp 1554483974
transform 1 0 1156 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_16
timestamp 1554483974
transform 1 0 1156 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_53
timestamp 1554483974
transform 1 0 1148 0 1 1515
box -2 -2 2 2
use M2_M1  M2_M1_56
timestamp 1554483974
transform 1 0 1132 0 1 1505
box -2 -2 2 2
use M3_M2  M3_M2_69
timestamp 1554483974
transform 1 0 1148 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_23
timestamp 1554483974
transform 1 0 1204 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_24
timestamp 1554483974
transform 1 0 1244 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_27
timestamp 1554483974
transform 1 0 1228 0 1 1555
box -3 -3 3 3
use M3_M2  M3_M2_42
timestamp 1554483974
transform 1 0 1228 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_17
timestamp 1554483974
transform 1 0 1220 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_18
timestamp 1554483974
transform 1 0 1228 0 1 1535
box -2 -2 2 2
use M3_M2  M3_M2_52
timestamp 1554483974
transform 1 0 1204 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_25
timestamp 1554483974
transform 1 0 1284 0 1 1565
box -3 -3 3 3
use M3_M2  M3_M2_43
timestamp 1554483974
transform 1 0 1276 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_41
timestamp 1554483974
transform 1 0 1244 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_70
timestamp 1554483974
transform 1 0 1244 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_19
timestamp 1554483974
transform 1 0 1292 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_42
timestamp 1554483974
transform 1 0 1316 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_44
timestamp 1554483974
transform 1 0 1364 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_20
timestamp 1554483974
transform 1 0 1364 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_54
timestamp 1554483974
transform 1 0 1356 0 1 1515
box -2 -2 2 2
use M3_M2  M3_M2_71
timestamp 1554483974
transform 1 0 1356 0 1 1505
box -3 -3 3 3
use M3_M2  M3_M2_45
timestamp 1554483974
transform 1 0 1388 0 1 1545
box -3 -3 3 3
use M2_M1  M2_M1_43
timestamp 1554483974
transform 1 0 1380 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_72
timestamp 1554483974
transform 1 0 1380 0 1 1505
box -3 -3 3 3
use M2_M1  M2_M1_44
timestamp 1554483974
transform 1 0 1412 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_28
timestamp 1554483974
transform 1 0 1436 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_21
timestamp 1554483974
transform 1 0 1436 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_22
timestamp 1554483974
transform 1 0 1452 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_23
timestamp 1554483974
transform 1 0 1540 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_45
timestamp 1554483974
transform 1 0 1460 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_46
timestamp 1554483974
transform 1 0 1500 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_53
timestamp 1554483974
transform 1 0 1540 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_29
timestamp 1554483974
transform 1 0 1564 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_47
timestamp 1554483974
transform 1 0 1564 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_24
timestamp 1554483974
transform 1 0 1660 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_48
timestamp 1554483974
transform 1 0 1636 0 1 1525
box -2 -2 2 2
use M3_M2  M3_M2_54
timestamp 1554483974
transform 1 0 1660 0 1 1525
box -3 -3 3 3
use M3_M2  M3_M2_30
timestamp 1554483974
transform 1 0 1700 0 1 1555
box -3 -3 3 3
use M2_M1  M2_M1_25
timestamp 1554483974
transform 1 0 1700 0 1 1535
box -2 -2 2 2
use M2_M1  M2_M1_49
timestamp 1554483974
transform 1 0 1692 0 1 1525
box -2 -2 2 2
use M2_M1  M2_M1_55
timestamp 1554483974
transform 1 0 1684 0 1 1515
box -2 -2 2 2
use UART_VIA1  UART_VIA1_1
timestamp 1554483974
transform 1 0 1801 0 1 1570
box -10 -3 10 3
use UART_VIA1  UART_VIA1_2
timestamp 1554483974
transform 1 0 24 0 1 1470
box -10 -3 10 3
use FILL  FILL_0
timestamp 1554483974
transform 1 0 72 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_0
timestamp 1554483974
transform -1 0 176 0 -1 1570
box -8 -3 104 105
use FILL  FILL_1
timestamp 1554483974
transform 1 0 176 0 -1 1570
box -8 -3 16 105
use FILL  FILL_2
timestamp 1554483974
transform 1 0 184 0 -1 1570
box -8 -3 16 105
use FILL  FILL_3
timestamp 1554483974
transform 1 0 192 0 -1 1570
box -8 -3 16 105
use FILL  FILL_4
timestamp 1554483974
transform 1 0 200 0 -1 1570
box -8 -3 16 105
use FILL  FILL_5
timestamp 1554483974
transform 1 0 208 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_1
timestamp 1554483974
transform 1 0 216 0 -1 1570
box -8 -3 104 105
use FILL  FILL_6
timestamp 1554483974
transform 1 0 312 0 -1 1570
box -8 -3 16 105
use FILL  FILL_7
timestamp 1554483974
transform 1 0 320 0 -1 1570
box -8 -3 16 105
use FILL  FILL_8
timestamp 1554483974
transform 1 0 328 0 -1 1570
box -8 -3 16 105
use FILL  FILL_9
timestamp 1554483974
transform 1 0 336 0 -1 1570
box -8 -3 16 105
use FILL  FILL_10
timestamp 1554483974
transform 1 0 344 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_0
timestamp 1554483974
transform 1 0 352 0 -1 1570
box -9 -3 26 105
use FILL  FILL_11
timestamp 1554483974
transform 1 0 368 0 -1 1570
box -8 -3 16 105
use FILL  FILL_12
timestamp 1554483974
transform 1 0 376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_13
timestamp 1554483974
transform 1 0 384 0 -1 1570
box -8 -3 16 105
use FILL  FILL_14
timestamp 1554483974
transform 1 0 392 0 -1 1570
box -8 -3 16 105
use FILL  FILL_15
timestamp 1554483974
transform 1 0 400 0 -1 1570
box -8 -3 16 105
use OR2X1  OR2X1_0
timestamp 1554483974
transform 1 0 408 0 -1 1570
box -8 -3 40 105
use OAI21X1  OAI21X1_0
timestamp 1554483974
transform 1 0 440 0 -1 1570
box -8 -3 34 105
use FILL  FILL_16
timestamp 1554483974
transform 1 0 472 0 -1 1570
box -8 -3 16 105
use FILL  FILL_17
timestamp 1554483974
transform 1 0 480 0 -1 1570
box -8 -3 16 105
use FILL  FILL_18
timestamp 1554483974
transform 1 0 488 0 -1 1570
box -8 -3 16 105
use FILL  FILL_19
timestamp 1554483974
transform 1 0 496 0 -1 1570
box -8 -3 16 105
use FILL  FILL_20
timestamp 1554483974
transform 1 0 504 0 -1 1570
box -8 -3 16 105
use FILL  FILL_21
timestamp 1554483974
transform 1 0 512 0 -1 1570
box -8 -3 16 105
use FILL  FILL_22
timestamp 1554483974
transform 1 0 520 0 -1 1570
box -8 -3 16 105
use FILL  FILL_23
timestamp 1554483974
transform 1 0 528 0 -1 1570
box -8 -3 16 105
use OAI21X1  OAI21X1_1
timestamp 1554483974
transform 1 0 536 0 -1 1570
box -8 -3 34 105
use FILL  FILL_24
timestamp 1554483974
transform 1 0 568 0 -1 1570
box -8 -3 16 105
use FILL  FILL_25
timestamp 1554483974
transform 1 0 576 0 -1 1570
box -8 -3 16 105
use FILL  FILL_26
timestamp 1554483974
transform 1 0 584 0 -1 1570
box -8 -3 16 105
use FILL  FILL_27
timestamp 1554483974
transform 1 0 592 0 -1 1570
box -8 -3 16 105
use FILL  FILL_28
timestamp 1554483974
transform 1 0 600 0 -1 1570
box -8 -3 16 105
use FILL  FILL_29
timestamp 1554483974
transform 1 0 608 0 -1 1570
box -8 -3 16 105
use FILL  FILL_30
timestamp 1554483974
transform 1 0 616 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_2
timestamp 1554483974
transform 1 0 624 0 -1 1570
box -8 -3 104 105
use FILL  FILL_31
timestamp 1554483974
transform 1 0 720 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_1
timestamp 1554483974
transform 1 0 728 0 -1 1570
box -9 -3 26 105
use FILL  FILL_32
timestamp 1554483974
transform 1 0 744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_33
timestamp 1554483974
transform 1 0 752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_34
timestamp 1554483974
transform 1 0 760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_35
timestamp 1554483974
transform 1 0 768 0 -1 1570
box -8 -3 16 105
use FILL  FILL_36
timestamp 1554483974
transform 1 0 776 0 -1 1570
box -8 -3 16 105
use FILL  FILL_37
timestamp 1554483974
transform 1 0 784 0 -1 1570
box -8 -3 16 105
use FILL  FILL_38
timestamp 1554483974
transform 1 0 792 0 -1 1570
box -8 -3 16 105
use INVX2  INVX2_2
timestamp 1554483974
transform 1 0 800 0 -1 1570
box -9 -3 26 105
use FILL  FILL_39
timestamp 1554483974
transform 1 0 816 0 -1 1570
box -8 -3 16 105
use OAI22X1  OAI22X1_0
timestamp 1554483974
transform -1 0 864 0 -1 1570
box -8 -3 46 105
use FILL  FILL_40
timestamp 1554483974
transform 1 0 864 0 -1 1570
box -8 -3 16 105
use FILL  FILL_41
timestamp 1554483974
transform 1 0 872 0 -1 1570
box -8 -3 16 105
use FILL  FILL_42
timestamp 1554483974
transform 1 0 880 0 -1 1570
box -8 -3 16 105
use FILL  FILL_43
timestamp 1554483974
transform 1 0 888 0 -1 1570
box -8 -3 16 105
use FILL  FILL_44
timestamp 1554483974
transform 1 0 896 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_3
timestamp 1554483974
transform -1 0 1000 0 -1 1570
box -8 -3 104 105
use FILL  FILL_45
timestamp 1554483974
transform 1 0 1000 0 -1 1570
box -8 -3 16 105
use FILL  FILL_46
timestamp 1554483974
transform 1 0 1008 0 -1 1570
box -8 -3 16 105
use FILL  FILL_47
timestamp 1554483974
transform 1 0 1016 0 -1 1570
box -8 -3 16 105
use NOR2X1  NOR2X1_0
timestamp 1554483974
transform 1 0 1024 0 -1 1570
box -8 -3 32 105
use FILL  FILL_48
timestamp 1554483974
transform 1 0 1048 0 -1 1570
box -8 -3 16 105
use FILL  FILL_49
timestamp 1554483974
transform 1 0 1056 0 -1 1570
box -8 -3 16 105
use FILL  FILL_50
timestamp 1554483974
transform 1 0 1064 0 -1 1570
box -8 -3 16 105
use FILL  FILL_51
timestamp 1554483974
transform 1 0 1072 0 -1 1570
box -8 -3 16 105
use FILL  FILL_52
timestamp 1554483974
transform 1 0 1080 0 -1 1570
box -8 -3 16 105
use FILL  FILL_53
timestamp 1554483974
transform 1 0 1088 0 -1 1570
box -8 -3 16 105
use FILL  FILL_54
timestamp 1554483974
transform 1 0 1096 0 -1 1570
box -8 -3 16 105
use FILL  FILL_55
timestamp 1554483974
transform 1 0 1104 0 -1 1570
box -8 -3 16 105
use FILL  FILL_56
timestamp 1554483974
transform 1 0 1112 0 -1 1570
box -8 -3 16 105
use NAND3X1  NAND3X1_0
timestamp 1554483974
transform -1 0 1152 0 -1 1570
box -8 -3 40 105
use FILL  FILL_57
timestamp 1554483974
transform 1 0 1152 0 -1 1570
box -8 -3 16 105
use FILL  FILL_58
timestamp 1554483974
transform 1 0 1160 0 -1 1570
box -8 -3 16 105
use XNOR2X1  XNOR2X1_0
timestamp 1554483974
transform -1 0 1224 0 -1 1570
box -8 -3 64 105
use XNOR2X1  XNOR2X1_1
timestamp 1554483974
transform -1 0 1280 0 -1 1570
box -8 -3 64 105
use FILL  FILL_59
timestamp 1554483974
transform 1 0 1280 0 -1 1570
box -8 -3 16 105
use FILL  FILL_60
timestamp 1554483974
transform 1 0 1288 0 -1 1570
box -8 -3 16 105
use FILL  FILL_61
timestamp 1554483974
transform 1 0 1296 0 -1 1570
box -8 -3 16 105
use FILL  FILL_62
timestamp 1554483974
transform 1 0 1304 0 -1 1570
box -8 -3 16 105
use FILL  FILL_63
timestamp 1554483974
transform 1 0 1312 0 -1 1570
box -8 -3 16 105
use LATCH  LATCH_0
timestamp 1554483974
transform -1 0 1376 0 -1 1570
box -8 -3 64 105
use FILL  FILL_64
timestamp 1554483974
transform 1 0 1376 0 -1 1570
box -8 -3 16 105
use FILL  FILL_65
timestamp 1554483974
transform 1 0 1384 0 -1 1570
box -8 -3 16 105
use AND2X2  AND2X2_0
timestamp 1554483974
transform -1 0 1424 0 -1 1570
box -8 -3 40 105
use FILL  FILL_66
timestamp 1554483974
transform 1 0 1424 0 -1 1570
box -8 -3 16 105
use FILL  FILL_67
timestamp 1554483974
transform 1 0 1432 0 -1 1570
box -8 -3 16 105
use FILL  FILL_68
timestamp 1554483974
transform 1 0 1440 0 -1 1570
box -8 -3 16 105
use FILL  FILL_69
timestamp 1554483974
transform 1 0 1448 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_4
timestamp 1554483974
transform -1 0 1552 0 -1 1570
box -8 -3 104 105
use FILL  FILL_70
timestamp 1554483974
transform 1 0 1552 0 -1 1570
box -8 -3 16 105
use FILL  FILL_71
timestamp 1554483974
transform 1 0 1560 0 -1 1570
box -8 -3 16 105
use FILL  FILL_72
timestamp 1554483974
transform 1 0 1568 0 -1 1570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_5
timestamp 1554483974
transform -1 0 1672 0 -1 1570
box -8 -3 104 105
use FILL  FILL_73
timestamp 1554483974
transform 1 0 1672 0 -1 1570
box -8 -3 16 105
use NAND2X1  NAND2X1_0
timestamp 1554483974
transform -1 0 1704 0 -1 1570
box -8 -3 32 105
use FILL  FILL_74
timestamp 1554483974
transform 1 0 1704 0 -1 1570
box -8 -3 16 105
use FILL  FILL_75
timestamp 1554483974
transform 1 0 1712 0 -1 1570
box -8 -3 16 105
use FILL  FILL_76
timestamp 1554483974
transform 1 0 1720 0 -1 1570
box -8 -3 16 105
use FILL  FILL_77
timestamp 1554483974
transform 1 0 1728 0 -1 1570
box -8 -3 16 105
use FILL  FILL_78
timestamp 1554483974
transform 1 0 1736 0 -1 1570
box -8 -3 16 105
use FILL  FILL_79
timestamp 1554483974
transform 1 0 1744 0 -1 1570
box -8 -3 16 105
use FILL  FILL_80
timestamp 1554483974
transform 1 0 1752 0 -1 1570
box -8 -3 16 105
use FILL  FILL_81
timestamp 1554483974
transform 1 0 1760 0 -1 1570
box -8 -3 16 105
use FILL  FILL_82
timestamp 1554483974
transform 1 0 1768 0 -1 1570
box -8 -3 16 105
use UART_VIA1  UART_VIA1_3
timestamp 1554483974
transform 1 0 1825 0 1 1470
box -10 -3 10 3
use M3_M2  M3_M2_92
timestamp 1554483974
transform 1 0 108 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_103
timestamp 1554483974
transform 1 0 108 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_68
timestamp 1554483974
transform 1 0 140 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_104
timestamp 1554483974
transform 1 0 164 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_122
timestamp 1554483974
transform 1 0 164 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_93
timestamp 1554483974
transform 1 0 180 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_69
timestamp 1554483974
transform 1 0 180 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_105
timestamp 1554483974
transform 1 0 188 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_104
timestamp 1554483974
transform 1 0 228 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_70
timestamp 1554483974
transform 1 0 244 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_71
timestamp 1554483974
transform 1 0 252 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_105
timestamp 1554483974
transform 1 0 244 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_94
timestamp 1554483974
transform 1 0 268 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_106
timestamp 1554483974
transform 1 0 276 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_107
timestamp 1554483974
transform 1 0 300 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_72
timestamp 1554483974
transform 1 0 316 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_106
timestamp 1554483974
transform 1 0 316 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_58
timestamp 1554483974
transform 1 0 332 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_108
timestamp 1554483974
transform 1 0 364 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_140
timestamp 1554483974
transform 1 0 356 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_109
timestamp 1554483974
transform 1 0 380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_123
timestamp 1554483974
transform 1 0 380 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_110
timestamp 1554483974
transform 1 0 420 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_73
timestamp 1554483974
transform 1 0 436 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_74
timestamp 1554483974
transform 1 0 452 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_107
timestamp 1554483974
transform 1 0 436 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_111
timestamp 1554483974
transform 1 0 444 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_112
timestamp 1554483974
transform 1 0 460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_124
timestamp 1554483974
transform 1 0 452 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_59
timestamp 1554483974
transform 1 0 476 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_60
timestamp 1554483974
transform 1 0 532 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_75
timestamp 1554483974
transform 1 0 524 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_113
timestamp 1554483974
transform 1 0 532 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_61
timestamp 1554483974
transform 1 0 548 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_76
timestamp 1554483974
transform 1 0 556 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_114
timestamp 1554483974
transform 1 0 548 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_62
timestamp 1554483974
transform 1 0 572 0 1 1425
box -2 -2 2 2
use M3_M2  M3_M2_95
timestamp 1554483974
transform 1 0 604 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_115
timestamp 1554483974
transform 1 0 604 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_108
timestamp 1554483974
transform 1 0 620 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_112
timestamp 1554483974
transform 1 0 612 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_75
timestamp 1554483974
transform 1 0 692 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_96
timestamp 1554483974
transform 1 0 708 0 1 1425
box -3 -3 3 3
use M2_M1  M2_M1_77
timestamp 1554483974
transform 1 0 692 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_78
timestamp 1554483974
transform 1 0 708 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_116
timestamp 1554483974
transform 1 0 700 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_76
timestamp 1554483974
transform 1 0 740 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_80
timestamp 1554483974
transform 1 0 732 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_97
timestamp 1554483974
transform 1 0 748 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_117
timestamp 1554483974
transform 1 0 748 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_79
timestamp 1554483974
transform 1 0 780 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_80
timestamp 1554483974
transform 1 0 804 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_118
timestamp 1554483974
transform 1 0 796 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_109
timestamp 1554483974
transform 1 0 804 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_119
timestamp 1554483974
transform 1 0 812 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_125
timestamp 1554483974
transform 1 0 796 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_77
timestamp 1554483974
transform 1 0 836 0 1 1455
box -3 -3 3 3
use M3_M2  M3_M2_84
timestamp 1554483974
transform 1 0 844 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_81
timestamp 1554483974
transform 1 0 836 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_113
timestamp 1554483974
transform 1 0 836 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_85
timestamp 1554483974
transform 1 0 876 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_98
timestamp 1554483974
transform 1 0 852 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_82
timestamp 1554483974
transform 1 0 876 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_83
timestamp 1554483974
transform 1 0 900 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_120
timestamp 1554483974
transform 1 0 852 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_121
timestamp 1554483974
transform 1 0 900 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_122
timestamp 1554483974
transform 1 0 908 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_114
timestamp 1554483974
transform 1 0 900 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_84
timestamp 1554483974
transform 1 0 924 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_115
timestamp 1554483974
transform 1 0 916 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_126
timestamp 1554483974
transform 1 0 916 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_99
timestamp 1554483974
transform 1 0 988 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_81
timestamp 1554483974
transform 1 0 1052 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_85
timestamp 1554483974
transform 1 0 1020 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_86
timestamp 1554483974
transform 1 0 1044 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_87
timestamp 1554483974
transform 1 0 1052 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_123
timestamp 1554483974
transform 1 0 964 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_127
timestamp 1554483974
transform 1 0 964 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_124
timestamp 1554483974
transform 1 0 1012 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_125
timestamp 1554483974
transform 1 0 1020 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_116
timestamp 1554483974
transform 1 0 1020 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_82
timestamp 1554483974
transform 1 0 1108 0 1 1445
box -3 -3 3 3
use M3_M2  M3_M2_86
timestamp 1554483974
transform 1 0 1108 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_100
timestamp 1554483974
transform 1 0 1092 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_83
timestamp 1554483974
transform 1 0 1148 0 1 1445
box -3 -3 3 3
use M2_M1  M2_M1_88
timestamp 1554483974
transform 1 0 1108 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_89
timestamp 1554483974
transform 1 0 1132 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_126
timestamp 1554483974
transform 1 0 1068 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_117
timestamp 1554483974
transform 1 0 1068 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_128
timestamp 1554483974
transform 1 0 1044 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_101
timestamp 1554483974
transform 1 0 1140 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_127
timestamp 1554483974
transform 1 0 1132 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_118
timestamp 1554483974
transform 1 0 1132 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_129
timestamp 1554483974
transform 1 0 1084 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_90
timestamp 1554483974
transform 1 0 1156 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_141
timestamp 1554483974
transform 1 0 1148 0 1 1395
box -2 -2 2 2
use M2_M1  M2_M1_142
timestamp 1554483974
transform 1 0 1164 0 1 1395
box -2 -2 2 2
use M3_M2  M3_M2_87
timestamp 1554483974
transform 1 0 1180 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_57
timestamp 1554483974
transform 1 0 1188 0 1 1435
box -2 -2 2 2
use M2_M1  M2_M1_63
timestamp 1554483974
transform 1 0 1260 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_91
timestamp 1554483974
transform 1 0 1228 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_128
timestamp 1554483974
transform 1 0 1212 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_64
timestamp 1554483974
transform 1 0 1316 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_92
timestamp 1554483974
transform 1 0 1284 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_129
timestamp 1554483974
transform 1 0 1268 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_102
timestamp 1554483974
transform 1 0 1316 0 1 1415
box -3 -3 3 3
use M3_M2  M3_M2_88
timestamp 1554483974
transform 1 0 1372 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_89
timestamp 1554483974
transform 1 0 1396 0 1 1435
box -3 -3 3 3
use M3_M2  M3_M2_90
timestamp 1554483974
transform 1 0 1412 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_65
timestamp 1554483974
transform 1 0 1372 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_93
timestamp 1554483974
transform 1 0 1340 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_130
timestamp 1554483974
transform 1 0 1324 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_119
timestamp 1554483974
transform 1 0 1284 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_91
timestamp 1554483974
transform 1 0 1444 0 1 1435
box -3 -3 3 3
use M2_M1  M2_M1_94
timestamp 1554483974
transform 1 0 1396 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_95
timestamp 1554483974
transform 1 0 1412 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_131
timestamp 1554483974
transform 1 0 1380 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_103
timestamp 1554483974
transform 1 0 1420 0 1 1415
box -3 -3 3 3
use M2_M1  M2_M1_96
timestamp 1554483974
transform 1 0 1428 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_97
timestamp 1554483974
transform 1 0 1444 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_132
timestamp 1554483974
transform 1 0 1420 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_120
timestamp 1554483974
transform 1 0 1420 0 1 1395
box -3 -3 3 3
use M2_M1  M2_M1_133
timestamp 1554483974
transform 1 0 1452 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_134
timestamp 1554483974
transform 1 0 1460 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_121
timestamp 1554483974
transform 1 0 1460 0 1 1395
box -3 -3 3 3
use M3_M2  M3_M2_130
timestamp 1554483974
transform 1 0 1452 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_66
timestamp 1554483974
transform 1 0 1492 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_98
timestamp 1554483974
transform 1 0 1516 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_135
timestamp 1554483974
transform 1 0 1500 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_99
timestamp 1554483974
transform 1 0 1532 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_136
timestamp 1554483974
transform 1 0 1524 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_131
timestamp 1554483974
transform 1 0 1532 0 1 1385
box -3 -3 3 3
use M2_M1  M2_M1_100
timestamp 1554483974
transform 1 0 1556 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_78
timestamp 1554483974
transform 1 0 1636 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_101
timestamp 1554483974
transform 1 0 1620 0 1 1415
box -2 -2 2 2
use M3_M2  M3_M2_110
timestamp 1554483974
transform 1 0 1620 0 1 1405
box -3 -3 3 3
use M2_M1  M2_M1_137
timestamp 1554483974
transform 1 0 1644 0 1 1405
box -2 -2 2 2
use M3_M2  M3_M2_132
timestamp 1554483974
transform 1 0 1628 0 1 1385
box -3 -3 3 3
use M3_M2  M3_M2_111
timestamp 1554483974
transform 1 0 1660 0 1 1405
box -3 -3 3 3
use M3_M2  M3_M2_79
timestamp 1554483974
transform 1 0 1700 0 1 1455
box -3 -3 3 3
use M2_M1  M2_M1_67
timestamp 1554483974
transform 1 0 1692 0 1 1425
box -2 -2 2 2
use M2_M1  M2_M1_102
timestamp 1554483974
transform 1 0 1676 0 1 1415
box -2 -2 2 2
use M2_M1  M2_M1_138
timestamp 1554483974
transform 1 0 1668 0 1 1405
box -2 -2 2 2
use M2_M1  M2_M1_139
timestamp 1554483974
transform 1 0 1700 0 1 1405
box -2 -2 2 2
use UART_VIA1  UART_VIA1_4
timestamp 1554483974
transform 1 0 48 0 1 1370
box -10 -3 10 3
use FILL  FILL_83
timestamp 1554483974
transform 1 0 72 0 1 1370
box -8 -3 16 105
use FILL  FILL_85
timestamp 1554483974
transform 1 0 80 0 1 1370
box -8 -3 16 105
use FILL  FILL_87
timestamp 1554483974
transform 1 0 88 0 1 1370
box -8 -3 16 105
use FILL  FILL_89
timestamp 1554483974
transform 1 0 96 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_3
timestamp 1554483974
transform 1 0 104 0 1 1370
box -9 -3 26 105
use FILL  FILL_91
timestamp 1554483974
transform 1 0 120 0 1 1370
box -8 -3 16 105
use FILL  FILL_95
timestamp 1554483974
transform 1 0 128 0 1 1370
box -8 -3 16 105
use FILL  FILL_97
timestamp 1554483974
transform 1 0 136 0 1 1370
box -8 -3 16 105
use FILL  FILL_99
timestamp 1554483974
transform 1 0 144 0 1 1370
box -8 -3 16 105
use FILL  FILL_101
timestamp 1554483974
transform 1 0 152 0 1 1370
box -8 -3 16 105
use FILL  FILL_103
timestamp 1554483974
transform 1 0 160 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_1
timestamp 1554483974
transform -1 0 208 0 1 1370
box -8 -3 46 105
use FILL  FILL_104
timestamp 1554483974
transform 1 0 208 0 1 1370
box -8 -3 16 105
use FILL  FILL_108
timestamp 1554483974
transform 1 0 216 0 1 1370
box -8 -3 16 105
use FILL  FILL_110
timestamp 1554483974
transform 1 0 224 0 1 1370
box -8 -3 16 105
use FILL  FILL_112
timestamp 1554483974
transform 1 0 232 0 1 1370
box -8 -3 16 105
use FILL  FILL_114
timestamp 1554483974
transform 1 0 240 0 1 1370
box -8 -3 16 105
use FILL  FILL_116
timestamp 1554483974
transform 1 0 248 0 1 1370
box -8 -3 16 105
use FILL  FILL_117
timestamp 1554483974
transform 1 0 256 0 1 1370
box -8 -3 16 105
use FILL  FILL_118
timestamp 1554483974
transform 1 0 264 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_2
timestamp 1554483974
transform 1 0 272 0 1 1370
box -8 -3 34 105
use FILL  FILL_119
timestamp 1554483974
transform 1 0 304 0 1 1370
box -8 -3 16 105
use FILL  FILL_125
timestamp 1554483974
transform 1 0 312 0 1 1370
box -8 -3 16 105
use FILL  FILL_126
timestamp 1554483974
transform 1 0 320 0 1 1370
box -8 -3 16 105
use FILL  FILL_127
timestamp 1554483974
transform 1 0 328 0 1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_1
timestamp 1554483974
transform -1 0 360 0 1 1370
box -8 -3 32 105
use FILL  FILL_128
timestamp 1554483974
transform 1 0 360 0 1 1370
box -8 -3 16 105
use FILL  FILL_131
timestamp 1554483974
transform 1 0 368 0 1 1370
box -8 -3 16 105
use FILL  FILL_133
timestamp 1554483974
transform 1 0 376 0 1 1370
box -8 -3 16 105
use FILL  FILL_135
timestamp 1554483974
transform 1 0 384 0 1 1370
box -8 -3 16 105
use FILL  FILL_137
timestamp 1554483974
transform 1 0 392 0 1 1370
box -8 -3 16 105
use FILL  FILL_139
timestamp 1554483974
transform 1 0 400 0 1 1370
box -8 -3 16 105
use FILL  FILL_141
timestamp 1554483974
transform 1 0 408 0 1 1370
box -8 -3 16 105
use FILL  FILL_143
timestamp 1554483974
transform 1 0 416 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_4
timestamp 1554483974
transform 1 0 424 0 1 1370
box -9 -3 26 105
use NAND2X1  NAND2X1_2
timestamp 1554483974
transform 1 0 440 0 1 1370
box -8 -3 32 105
use FILL  FILL_145
timestamp 1554483974
transform 1 0 464 0 1 1370
box -8 -3 16 105
use FILL  FILL_149
timestamp 1554483974
transform 1 0 472 0 1 1370
box -8 -3 16 105
use FILL  FILL_151
timestamp 1554483974
transform 1 0 480 0 1 1370
box -8 -3 16 105
use FILL  FILL_153
timestamp 1554483974
transform 1 0 488 0 1 1370
box -8 -3 16 105
use FILL  FILL_155
timestamp 1554483974
transform 1 0 496 0 1 1370
box -8 -3 16 105
use FILL  FILL_157
timestamp 1554483974
transform 1 0 504 0 1 1370
box -8 -3 16 105
use FILL  FILL_159
timestamp 1554483974
transform 1 0 512 0 1 1370
box -8 -3 16 105
use FILL  FILL_161
timestamp 1554483974
transform 1 0 520 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_3
timestamp 1554483974
transform 1 0 528 0 1 1370
box -8 -3 32 105
use NAND2X1  NAND2X1_4
timestamp 1554483974
transform 1 0 552 0 1 1370
box -8 -3 32 105
use FILL  FILL_163
timestamp 1554483974
transform 1 0 576 0 1 1370
box -8 -3 16 105
use FILL  FILL_167
timestamp 1554483974
transform 1 0 584 0 1 1370
box -8 -3 16 105
use FILL  FILL_169
timestamp 1554483974
transform 1 0 592 0 1 1370
box -8 -3 16 105
use FILL  FILL_171
timestamp 1554483974
transform 1 0 600 0 1 1370
box -8 -3 16 105
use FILL  FILL_172
timestamp 1554483974
transform 1 0 608 0 1 1370
box -8 -3 16 105
use FILL  FILL_173
timestamp 1554483974
transform 1 0 616 0 1 1370
box -8 -3 16 105
use FILL  FILL_174
timestamp 1554483974
transform 1 0 624 0 1 1370
box -8 -3 16 105
use FILL  FILL_175
timestamp 1554483974
transform 1 0 632 0 1 1370
box -8 -3 16 105
use INVX2  INVX2_5
timestamp 1554483974
transform 1 0 640 0 1 1370
box -9 -3 26 105
use FILL  FILL_176
timestamp 1554483974
transform 1 0 656 0 1 1370
box -8 -3 16 105
use FILL  FILL_177
timestamp 1554483974
transform 1 0 664 0 1 1370
box -8 -3 16 105
use FILL  FILL_178
timestamp 1554483974
transform 1 0 672 0 1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_2
timestamp 1554483974
transform -1 0 720 0 1 1370
box -8 -3 46 105
use FILL  FILL_179
timestamp 1554483974
transform 1 0 720 0 1 1370
box -8 -3 16 105
use FILL  FILL_189
timestamp 1554483974
transform 1 0 728 0 1 1370
box -8 -3 16 105
use FILL  FILL_190
timestamp 1554483974
transform 1 0 736 0 1 1370
box -8 -3 16 105
use FILL  FILL_191
timestamp 1554483974
transform 1 0 744 0 1 1370
box -8 -3 16 105
use FILL  FILL_192
timestamp 1554483974
transform 1 0 752 0 1 1370
box -8 -3 16 105
use FILL  FILL_193
timestamp 1554483974
transform 1 0 760 0 1 1370
box -8 -3 16 105
use FILL  FILL_194
timestamp 1554483974
transform 1 0 768 0 1 1370
box -8 -3 16 105
use FILL  FILL_195
timestamp 1554483974
transform 1 0 776 0 1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_1
timestamp 1554483974
transform -1 0 824 0 1 1370
box -8 -3 46 105
use FILL  FILL_196
timestamp 1554483974
transform 1 0 824 0 1 1370
box -8 -3 16 105
use FILL  FILL_197
timestamp 1554483974
transform 1 0 832 0 1 1370
box -8 -3 16 105
use FILL  FILL_198
timestamp 1554483974
transform 1 0 840 0 1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_0
timestamp 1554483974
transform 1 0 848 0 1 1370
box -8 -3 64 105
use FILL  FILL_199
timestamp 1554483974
transform 1 0 904 0 1 1370
box -8 -3 16 105
use FILL  FILL_200
timestamp 1554483974
transform 1 0 912 0 1 1370
box -8 -3 16 105
use FILL  FILL_207
timestamp 1554483974
transform 1 0 920 0 1 1370
box -8 -3 16 105
use FILL  FILL_209
timestamp 1554483974
transform 1 0 928 0 1 1370
box -8 -3 16 105
use FILL  FILL_211
timestamp 1554483974
transform 1 0 936 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_133
timestamp 1554483974
transform 1 0 956 0 1 1375
box -3 -3 3 3
use INVX2  INVX2_8
timestamp 1554483974
transform 1 0 944 0 1 1370
box -9 -3 26 105
use M3_M2  M3_M2_134
timestamp 1554483974
transform 1 0 988 0 1 1375
box -3 -3 3 3
use XOR2X1  XOR2X1_2
timestamp 1554483974
transform 1 0 960 0 1 1370
box -8 -3 64 105
use XOR2X1  XOR2X1_3
timestamp 1554483974
transform 1 0 1016 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_135
timestamp 1554483974
transform 1 0 1092 0 1 1375
box -3 -3 3 3
use XNOR2X1  XNOR2X1_2
timestamp 1554483974
transform 1 0 1072 0 1 1370
box -8 -3 64 105
use NOR2X1  NOR2X1_3
timestamp 1554483974
transform -1 0 1152 0 1 1370
box -8 -3 32 105
use FILL  FILL_212
timestamp 1554483974
transform 1 0 1152 0 1 1370
box -8 -3 16 105
use FILL  FILL_213
timestamp 1554483974
transform 1 0 1160 0 1 1370
box -8 -3 16 105
use M3_M2  M3_M2_136
timestamp 1554483974
transform 1 0 1180 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_137
timestamp 1554483974
transform 1 0 1212 0 1 1375
box -3 -3 3 3
use LATCH  LATCH_1
timestamp 1554483974
transform -1 0 1224 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_138
timestamp 1554483974
transform 1 0 1252 0 1 1375
box -3 -3 3 3
use M3_M2  M3_M2_139
timestamp 1554483974
transform 1 0 1268 0 1 1375
box -3 -3 3 3
use LATCH  LATCH_2
timestamp 1554483974
transform -1 0 1280 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_140
timestamp 1554483974
transform 1 0 1316 0 1 1375
box -3 -3 3 3
use LATCH  LATCH_3
timestamp 1554483974
transform -1 0 1336 0 1 1370
box -8 -3 64 105
use M3_M2  M3_M2_141
timestamp 1554483974
transform 1 0 1380 0 1 1375
box -3 -3 3 3
use LATCH  LATCH_4
timestamp 1554483974
transform -1 0 1392 0 1 1370
box -8 -3 64 105
use AND2X2  AND2X2_1
timestamp 1554483974
transform -1 0 1424 0 1 1370
box -8 -3 40 105
use AND2X2  AND2X2_2
timestamp 1554483974
transform -1 0 1456 0 1 1370
box -8 -3 40 105
use FILL  FILL_214
timestamp 1554483974
transform 1 0 1456 0 1 1370
box -8 -3 16 105
use FILL  FILL_242
timestamp 1554483974
transform 1 0 1464 0 1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_5
timestamp 1554483974
transform 1 0 1472 0 1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_5
timestamp 1554483974
transform -1 0 1528 0 1 1370
box -8 -3 34 105
use FILL  FILL_244
timestamp 1554483974
transform 1 0 1528 0 1 1370
box -8 -3 16 105
use FILL  FILL_245
timestamp 1554483974
transform 1 0 1536 0 1 1370
box -8 -3 16 105
use FILL  FILL_246
timestamp 1554483974
transform 1 0 1544 0 1 1370
box -8 -3 16 105
use FILL  FILL_247
timestamp 1554483974
transform 1 0 1552 0 1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_6
timestamp 1554483974
transform -1 0 1656 0 1 1370
box -8 -3 104 105
use FILL  FILL_248
timestamp 1554483974
transform 1 0 1656 0 1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_6
timestamp 1554483974
transform 1 0 1664 0 1 1370
box -8 -3 34 105
use FILL  FILL_249
timestamp 1554483974
transform 1 0 1696 0 1 1370
box -8 -3 16 105
use FILL  FILL_257
timestamp 1554483974
transform 1 0 1704 0 1 1370
box -8 -3 16 105
use FILL  FILL_259
timestamp 1554483974
transform 1 0 1712 0 1 1370
box -8 -3 16 105
use FILL  FILL_261
timestamp 1554483974
transform 1 0 1720 0 1 1370
box -8 -3 16 105
use FILL  FILL_263
timestamp 1554483974
transform 1 0 1728 0 1 1370
box -8 -3 16 105
use FILL  FILL_265
timestamp 1554483974
transform 1 0 1736 0 1 1370
box -8 -3 16 105
use FILL  FILL_267
timestamp 1554483974
transform 1 0 1744 0 1 1370
box -8 -3 16 105
use FILL  FILL_269
timestamp 1554483974
transform 1 0 1752 0 1 1370
box -8 -3 16 105
use FILL  FILL_271
timestamp 1554483974
transform 1 0 1760 0 1 1370
box -8 -3 16 105
use FILL  FILL_273
timestamp 1554483974
transform 1 0 1768 0 1 1370
box -8 -3 16 105
use UART_VIA1  UART_VIA1_5
timestamp 1554483974
transform 1 0 1801 0 1 1370
box -10 -3 10 3
use M3_M2  M3_M2_161
timestamp 1554483974
transform 1 0 140 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_211
timestamp 1554483974
transform 1 0 140 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_142
timestamp 1554483974
transform 1 0 156 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_179
timestamp 1554483974
transform 1 0 172 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_180
timestamp 1554483974
transform 1 0 172 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_222
timestamp 1554483974
transform 1 0 180 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_199
timestamp 1554483974
transform 1 0 180 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_143
timestamp 1554483974
transform 1 0 204 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_212
timestamp 1554483974
transform 1 0 196 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_200
timestamp 1554483974
transform 1 0 220 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_146
timestamp 1554483974
transform 1 0 244 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_181
timestamp 1554483974
transform 1 0 244 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_144
timestamp 1554483974
transform 1 0 284 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_180
timestamp 1554483974
transform 1 0 284 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_147
timestamp 1554483974
transform 1 0 316 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_162
timestamp 1554483974
transform 1 0 348 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_148
timestamp 1554483974
transform 1 0 348 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_181
timestamp 1554483974
transform 1 0 324 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_182
timestamp 1554483974
transform 1 0 340 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_183
timestamp 1554483974
transform 1 0 364 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_145
timestamp 1554483974
transform 1 0 404 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_143
timestamp 1554483974
transform 1 0 396 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_144
timestamp 1554483974
transform 1 0 436 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_149
timestamp 1554483974
transform 1 0 444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_184
timestamp 1554483974
transform 1 0 452 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_150
timestamp 1554483974
transform 1 0 468 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_189
timestamp 1554483974
transform 1 0 476 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_151
timestamp 1554483974
transform 1 0 516 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_152
timestamp 1554483974
transform 1 0 532 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_185
timestamp 1554483974
transform 1 0 524 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_172
timestamp 1554483974
transform 1 0 548 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_213
timestamp 1554483974
transform 1 0 556 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_146
timestamp 1554483974
transform 1 0 572 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_214
timestamp 1554483974
transform 1 0 588 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_163
timestamp 1554483974
transform 1 0 604 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_153
timestamp 1554483974
transform 1 0 604 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_154
timestamp 1554483974
transform 1 0 612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_155
timestamp 1554483974
transform 1 0 628 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_173
timestamp 1554483974
transform 1 0 636 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_147
timestamp 1554483974
transform 1 0 652 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_156
timestamp 1554483974
transform 1 0 652 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_186
timestamp 1554483974
transform 1 0 620 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_187
timestamp 1554483974
transform 1 0 636 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_188
timestamp 1554483974
transform 1 0 644 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_182
timestamp 1554483974
transform 1 0 644 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_189
timestamp 1554483974
transform 1 0 660 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_190
timestamp 1554483974
transform 1 0 660 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_148
timestamp 1554483974
transform 1 0 700 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_157
timestamp 1554483974
transform 1 0 700 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_164
timestamp 1554483974
transform 1 0 764 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_158
timestamp 1554483974
transform 1 0 756 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_159
timestamp 1554483974
transform 1 0 764 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_174
timestamp 1554483974
transform 1 0 772 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_190
timestamp 1554483974
transform 1 0 724 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_191
timestamp 1554483974
transform 1 0 732 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_192
timestamp 1554483974
transform 1 0 748 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_193
timestamp 1554483974
transform 1 0 764 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_191
timestamp 1554483974
transform 1 0 716 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_183
timestamp 1554483974
transform 1 0 748 0 1 1315
box -3 -3 3 3
use M3_M2  M3_M2_192
timestamp 1554483974
transform 1 0 764 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_194
timestamp 1554483974
transform 1 0 788 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_193
timestamp 1554483974
transform 1 0 780 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_149
timestamp 1554483974
transform 1 0 812 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_165
timestamp 1554483974
transform 1 0 820 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_157
timestamp 1554483974
transform 1 0 836 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_158
timestamp 1554483974
transform 1 0 852 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_175
timestamp 1554483974
transform 1 0 828 0 1 1335
box -3 -3 3 3
use M3_M2  M3_M2_166
timestamp 1554483974
transform 1 0 860 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_176
timestamp 1554483974
transform 1 0 852 0 1 1335
box -3 -3 3 3
use M2_M1  M2_M1_160
timestamp 1554483974
transform 1 0 860 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_195
timestamp 1554483974
transform 1 0 844 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_196
timestamp 1554483974
transform 1 0 860 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_215
timestamp 1554483974
transform 1 0 828 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_216
timestamp 1554483974
transform 1 0 852 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_223
timestamp 1554483974
transform 1 0 852 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_159
timestamp 1554483974
transform 1 0 908 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_201
timestamp 1554483974
transform 1 0 852 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_202
timestamp 1554483974
transform 1 0 884 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_150
timestamp 1554483974
transform 1 0 932 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_167
timestamp 1554483974
transform 1 0 932 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_161
timestamp 1554483974
transform 1 0 924 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_162
timestamp 1554483974
transform 1 0 932 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_160
timestamp 1554483974
transform 1 0 948 0 1 1355
box -3 -3 3 3
use M3_M2  M3_M2_177
timestamp 1554483974
transform 1 0 964 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_163
timestamp 1554483974
transform 1 0 1004 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_184
timestamp 1554483974
transform 1 0 1004 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_145
timestamp 1554483974
transform 1 0 1036 0 1 1345
box -2 -2 2 2
use M2_M1  M2_M1_164
timestamp 1554483974
transform 1 0 1052 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_203
timestamp 1554483974
transform 1 0 1052 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_185
timestamp 1554483974
transform 1 0 1068 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_197
timestamp 1554483974
transform 1 0 1092 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_217
timestamp 1554483974
transform 1 0 1076 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_218
timestamp 1554483974
transform 1 0 1100 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_224
timestamp 1554483974
transform 1 0 1084 0 1 1305
box -2 -2 2 2
use M3_M2  M3_M2_204
timestamp 1554483974
transform 1 0 1084 0 1 1295
box -3 -3 3 3
use M2_M1  M2_M1_165
timestamp 1554483974
transform 1 0 1156 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_166
timestamp 1554483974
transform 1 0 1188 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_167
timestamp 1554483974
transform 1 0 1204 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_198
timestamp 1554483974
transform 1 0 1164 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_199
timestamp 1554483974
transform 1 0 1180 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_200
timestamp 1554483974
transform 1 0 1196 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_194
timestamp 1554483974
transform 1 0 1164 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_195
timestamp 1554483974
transform 1 0 1196 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_201
timestamp 1554483974
transform 1 0 1220 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_151
timestamp 1554483974
transform 1 0 1268 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_202
timestamp 1554483974
transform 1 0 1244 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_203
timestamp 1554483974
transform 1 0 1260 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_196
timestamp 1554483974
transform 1 0 1244 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_205
timestamp 1554483974
transform 1 0 1244 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_152
timestamp 1554483974
transform 1 0 1300 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_168
timestamp 1554483974
transform 1 0 1316 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_204
timestamp 1554483974
transform 1 0 1276 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_186
timestamp 1554483974
transform 1 0 1276 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_219
timestamp 1554483974
transform 1 0 1308 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_197
timestamp 1554483974
transform 1 0 1308 0 1 1305
box -3 -3 3 3
use M2_M1  M2_M1_205
timestamp 1554483974
transform 1 0 1332 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_198
timestamp 1554483974
transform 1 0 1332 0 1 1305
box -3 -3 3 3
use M3_M2  M3_M2_206
timestamp 1554483974
transform 1 0 1356 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_153
timestamp 1554483974
transform 1 0 1420 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_168
timestamp 1554483974
transform 1 0 1404 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_169
timestamp 1554483974
transform 1 0 1404 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_170
timestamp 1554483974
transform 1 0 1412 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_206
timestamp 1554483974
transform 1 0 1396 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_207
timestamp 1554483974
transform 1 0 1412 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_207
timestamp 1554483974
transform 1 0 1396 0 1 1295
box -3 -3 3 3
use M3_M2  M3_M2_169
timestamp 1554483974
transform 1 0 1444 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_171
timestamp 1554483974
transform 1 0 1436 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_187
timestamp 1554483974
transform 1 0 1436 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_172
timestamp 1554483974
transform 1 0 1444 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_173
timestamp 1554483974
transform 1 0 1476 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_174
timestamp 1554483974
transform 1 0 1492 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_208
timestamp 1554483974
transform 1 0 1508 0 1 1325
box -2 -2 2 2
use M2_M1  M2_M1_220
timestamp 1554483974
transform 1 0 1508 0 1 1315
box -2 -2 2 2
use M3_M2  M3_M2_154
timestamp 1554483974
transform 1 0 1524 0 1 1365
box -3 -3 3 3
use M3_M2  M3_M2_170
timestamp 1554483974
transform 1 0 1612 0 1 1345
box -3 -3 3 3
use M2_M1  M2_M1_175
timestamp 1554483974
transform 1 0 1612 0 1 1335
box -2 -2 2 2
use M2_M1  M2_M1_209
timestamp 1554483974
transform 1 0 1564 0 1 1325
box -2 -2 2 2
use M3_M2  M3_M2_188
timestamp 1554483974
transform 1 0 1564 0 1 1315
box -3 -3 3 3
use M2_M1  M2_M1_176
timestamp 1554483974
transform 1 0 1628 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_171
timestamp 1554483974
transform 1 0 1644 0 1 1345
box -3 -3 3 3
use M3_M2  M3_M2_155
timestamp 1554483974
transform 1 0 1668 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_177
timestamp 1554483974
transform 1 0 1660 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_156
timestamp 1554483974
transform 1 0 1692 0 1 1365
box -3 -3 3 3
use M2_M1  M2_M1_178
timestamp 1554483974
transform 1 0 1692 0 1 1335
box -2 -2 2 2
use M3_M2  M3_M2_178
timestamp 1554483974
transform 1 0 1660 0 1 1325
box -3 -3 3 3
use M3_M2  M3_M2_179
timestamp 1554483974
transform 1 0 1684 0 1 1325
box -3 -3 3 3
use M2_M1  M2_M1_221
timestamp 1554483974
transform 1 0 1660 0 1 1315
box -2 -2 2 2
use M2_M1  M2_M1_210
timestamp 1554483974
transform 1 0 1716 0 1 1325
box -2 -2 2 2
use UART_VIA1  UART_VIA1_6
timestamp 1554483974
transform 1 0 24 0 1 1270
box -10 -3 10 3
use FILL  FILL_84
timestamp 1554483974
transform 1 0 72 0 -1 1370
box -8 -3 16 105
use FILL  FILL_86
timestamp 1554483974
transform 1 0 80 0 -1 1370
box -8 -3 16 105
use FILL  FILL_88
timestamp 1554483974
transform 1 0 88 0 -1 1370
box -8 -3 16 105
use FILL  FILL_90
timestamp 1554483974
transform 1 0 96 0 -1 1370
box -8 -3 16 105
use FILL  FILL_92
timestamp 1554483974
transform 1 0 104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_93
timestamp 1554483974
transform 1 0 112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_94
timestamp 1554483974
transform 1 0 120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_96
timestamp 1554483974
transform 1 0 128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_98
timestamp 1554483974
transform 1 0 136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_100
timestamp 1554483974
transform 1 0 144 0 -1 1370
box -8 -3 16 105
use FILL  FILL_102
timestamp 1554483974
transform 1 0 152 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_1
timestamp 1554483974
transform 1 0 160 0 -1 1370
box -8 -3 40 105
use FILL  FILL_105
timestamp 1554483974
transform 1 0 192 0 -1 1370
box -8 -3 16 105
use FILL  FILL_106
timestamp 1554483974
transform 1 0 200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_107
timestamp 1554483974
transform 1 0 208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_109
timestamp 1554483974
transform 1 0 216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_111
timestamp 1554483974
transform 1 0 224 0 -1 1370
box -8 -3 16 105
use FILL  FILL_113
timestamp 1554483974
transform 1 0 232 0 -1 1370
box -8 -3 16 105
use FILL  FILL_115
timestamp 1554483974
transform 1 0 240 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_1
timestamp 1554483974
transform 1 0 248 0 -1 1370
box -8 -3 32 105
use FILL  FILL_120
timestamp 1554483974
transform 1 0 272 0 -1 1370
box -8 -3 16 105
use FILL  FILL_121
timestamp 1554483974
transform 1 0 280 0 -1 1370
box -8 -3 16 105
use FILL  FILL_122
timestamp 1554483974
transform 1 0 288 0 -1 1370
box -8 -3 16 105
use FILL  FILL_123
timestamp 1554483974
transform 1 0 296 0 -1 1370
box -8 -3 16 105
use FILL  FILL_124
timestamp 1554483974
transform 1 0 304 0 -1 1370
box -8 -3 16 105
use FILL  FILL_129
timestamp 1554483974
transform 1 0 312 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_0
timestamp 1554483974
transform -1 0 360 0 -1 1370
box -8 -3 46 105
use FILL  FILL_130
timestamp 1554483974
transform 1 0 360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_132
timestamp 1554483974
transform 1 0 368 0 -1 1370
box -8 -3 16 105
use FILL  FILL_134
timestamp 1554483974
transform 1 0 376 0 -1 1370
box -8 -3 16 105
use FILL  FILL_136
timestamp 1554483974
transform 1 0 384 0 -1 1370
box -8 -3 16 105
use FILL  FILL_138
timestamp 1554483974
transform 1 0 392 0 -1 1370
box -8 -3 16 105
use FILL  FILL_140
timestamp 1554483974
transform 1 0 400 0 -1 1370
box -8 -3 16 105
use FILL  FILL_142
timestamp 1554483974
transform 1 0 408 0 -1 1370
box -8 -3 16 105
use FILL  FILL_144
timestamp 1554483974
transform 1 0 416 0 -1 1370
box -8 -3 16 105
use FILL  FILL_146
timestamp 1554483974
transform 1 0 424 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_2
timestamp 1554483974
transform 1 0 432 0 -1 1370
box -8 -3 32 105
use FILL  FILL_147
timestamp 1554483974
transform 1 0 456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_148
timestamp 1554483974
transform 1 0 464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_150
timestamp 1554483974
transform 1 0 472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_152
timestamp 1554483974
transform 1 0 480 0 -1 1370
box -8 -3 16 105
use FILL  FILL_154
timestamp 1554483974
transform 1 0 488 0 -1 1370
box -8 -3 16 105
use FILL  FILL_156
timestamp 1554483974
transform 1 0 496 0 -1 1370
box -8 -3 16 105
use FILL  FILL_158
timestamp 1554483974
transform 1 0 504 0 -1 1370
box -8 -3 16 105
use FILL  FILL_160
timestamp 1554483974
transform 1 0 512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_162
timestamp 1554483974
transform 1 0 520 0 -1 1370
box -8 -3 16 105
use OAI21X1  OAI21X1_3
timestamp 1554483974
transform 1 0 528 0 -1 1370
box -8 -3 34 105
use FILL  FILL_164
timestamp 1554483974
transform 1 0 560 0 -1 1370
box -8 -3 16 105
use FILL  FILL_165
timestamp 1554483974
transform 1 0 568 0 -1 1370
box -8 -3 16 105
use FILL  FILL_166
timestamp 1554483974
transform 1 0 576 0 -1 1370
box -8 -3 16 105
use FILL  FILL_168
timestamp 1554483974
transform 1 0 584 0 -1 1370
box -8 -3 16 105
use FILL  FILL_170
timestamp 1554483974
transform 1 0 592 0 -1 1370
box -8 -3 16 105
use FILL  FILL_180
timestamp 1554483974
transform 1 0 600 0 -1 1370
box -8 -3 16 105
use OAI22X1  OAI22X1_3
timestamp 1554483974
transform -1 0 648 0 -1 1370
box -8 -3 46 105
use FILL  FILL_181
timestamp 1554483974
transform 1 0 648 0 -1 1370
box -8 -3 16 105
use INVX2  INVX2_6
timestamp 1554483974
transform 1 0 656 0 -1 1370
box -9 -3 26 105
use FILL  FILL_182
timestamp 1554483974
transform 1 0 672 0 -1 1370
box -8 -3 16 105
use FILL  FILL_183
timestamp 1554483974
transform 1 0 680 0 -1 1370
box -8 -3 16 105
use FILL  FILL_184
timestamp 1554483974
transform 1 0 688 0 -1 1370
box -8 -3 16 105
use FILL  FILL_185
timestamp 1554483974
transform 1 0 696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_186
timestamp 1554483974
transform 1 0 704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_187
timestamp 1554483974
transform 1 0 712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_188
timestamp 1554483974
transform 1 0 720 0 -1 1370
box -8 -3 16 105
use AOI22X1  AOI22X1_2
timestamp 1554483974
transform 1 0 728 0 -1 1370
box -8 -3 46 105
use INVX2  INVX2_7
timestamp 1554483974
transform 1 0 768 0 -1 1370
box -9 -3 26 105
use FILL  FILL_201
timestamp 1554483974
transform 1 0 784 0 -1 1370
box -8 -3 16 105
use FILL  FILL_202
timestamp 1554483974
transform 1 0 792 0 -1 1370
box -8 -3 16 105
use FILL  FILL_203
timestamp 1554483974
transform 1 0 800 0 -1 1370
box -8 -3 16 105
use FILL  FILL_204
timestamp 1554483974
transform 1 0 808 0 -1 1370
box -8 -3 16 105
use FILL  FILL_205
timestamp 1554483974
transform 1 0 816 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_2
timestamp 1554483974
transform -1 0 856 0 -1 1370
box -8 -3 40 105
use XOR2X1  XOR2X1_1
timestamp 1554483974
transform -1 0 912 0 -1 1370
box -8 -3 64 105
use FILL  FILL_206
timestamp 1554483974
transform 1 0 912 0 -1 1370
box -8 -3 16 105
use FILL  FILL_208
timestamp 1554483974
transform 1 0 920 0 -1 1370
box -8 -3 16 105
use FILL  FILL_210
timestamp 1554483974
transform 1 0 928 0 -1 1370
box -8 -3 16 105
use XOR2X1  XOR2X1_4
timestamp 1554483974
transform 1 0 936 0 -1 1370
box -8 -3 64 105
use FILL  FILL_215
timestamp 1554483974
transform 1 0 992 0 -1 1370
box -8 -3 16 105
use FILL  FILL_216
timestamp 1554483974
transform 1 0 1000 0 -1 1370
box -8 -3 16 105
use NOR2X1  NOR2X1_4
timestamp 1554483974
transform -1 0 1032 0 -1 1370
box -8 -3 32 105
use FILL  FILL_217
timestamp 1554483974
transform 1 0 1032 0 -1 1370
box -8 -3 16 105
use FILL  FILL_218
timestamp 1554483974
transform 1 0 1040 0 -1 1370
box -8 -3 16 105
use FILL  FILL_219
timestamp 1554483974
transform 1 0 1048 0 -1 1370
box -8 -3 16 105
use FILL  FILL_220
timestamp 1554483974
transform 1 0 1056 0 -1 1370
box -8 -3 16 105
use FILL  FILL_221
timestamp 1554483974
transform 1 0 1064 0 -1 1370
box -8 -3 16 105
use NAND3X1  NAND3X1_3
timestamp 1554483974
transform -1 0 1104 0 -1 1370
box -8 -3 40 105
use FILL  FILL_222
timestamp 1554483974
transform 1 0 1104 0 -1 1370
box -8 -3 16 105
use FILL  FILL_223
timestamp 1554483974
transform 1 0 1112 0 -1 1370
box -8 -3 16 105
use FILL  FILL_224
timestamp 1554483974
transform 1 0 1120 0 -1 1370
box -8 -3 16 105
use FILL  FILL_225
timestamp 1554483974
transform 1 0 1128 0 -1 1370
box -8 -3 16 105
use FILL  FILL_226
timestamp 1554483974
transform 1 0 1136 0 -1 1370
box -8 -3 16 105
use FILL  FILL_227
timestamp 1554483974
transform 1 0 1144 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_3
timestamp 1554483974
transform 1 0 1152 0 -1 1370
box -8 -3 40 105
use INVX2  INVX2_9
timestamp 1554483974
transform 1 0 1184 0 -1 1370
box -9 -3 26 105
use FILL  FILL_228
timestamp 1554483974
transform 1 0 1200 0 -1 1370
box -8 -3 16 105
use FILL  FILL_229
timestamp 1554483974
transform 1 0 1208 0 -1 1370
box -8 -3 16 105
use FILL  FILL_230
timestamp 1554483974
transform 1 0 1216 0 -1 1370
box -8 -3 16 105
use FILL  FILL_231
timestamp 1554483974
transform 1 0 1224 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_4
timestamp 1554483974
transform 1 0 1232 0 -1 1370
box -8 -3 40 105
use FILL  FILL_232
timestamp 1554483974
transform 1 0 1264 0 -1 1370
box -8 -3 16 105
use LATCH  LATCH_5
timestamp 1554483974
transform -1 0 1328 0 -1 1370
box -8 -3 64 105
use FILL  FILL_233
timestamp 1554483974
transform 1 0 1328 0 -1 1370
box -8 -3 16 105
use FILL  FILL_234
timestamp 1554483974
transform 1 0 1336 0 -1 1370
box -8 -3 16 105
use FILL  FILL_235
timestamp 1554483974
transform 1 0 1344 0 -1 1370
box -8 -3 16 105
use FILL  FILL_236
timestamp 1554483974
transform 1 0 1352 0 -1 1370
box -8 -3 16 105
use FILL  FILL_237
timestamp 1554483974
transform 1 0 1360 0 -1 1370
box -8 -3 16 105
use FILL  FILL_238
timestamp 1554483974
transform 1 0 1368 0 -1 1370
box -8 -3 16 105
use AND2X2  AND2X2_5
timestamp 1554483974
transform -1 0 1408 0 -1 1370
box -8 -3 40 105
use OAI21X1  OAI21X1_4
timestamp 1554483974
transform 1 0 1408 0 -1 1370
box -8 -3 34 105
use FILL  FILL_239
timestamp 1554483974
transform 1 0 1440 0 -1 1370
box -8 -3 16 105
use FILL  FILL_240
timestamp 1554483974
transform 1 0 1448 0 -1 1370
box -8 -3 16 105
use FILL  FILL_241
timestamp 1554483974
transform 1 0 1456 0 -1 1370
box -8 -3 16 105
use FILL  FILL_243
timestamp 1554483974
transform 1 0 1464 0 -1 1370
box -8 -3 16 105
use FILL  FILL_250
timestamp 1554483974
transform 1 0 1472 0 -1 1370
box -8 -3 16 105
use FILL  FILL_251
timestamp 1554483974
transform 1 0 1480 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_6
timestamp 1554483974
transform 1 0 1488 0 -1 1370
box -8 -3 32 105
use FILL  FILL_252
timestamp 1554483974
transform 1 0 1512 0 -1 1370
box -8 -3 16 105
use FILL  FILL_253
timestamp 1554483974
transform 1 0 1520 0 -1 1370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_7
timestamp 1554483974
transform -1 0 1624 0 -1 1370
box -8 -3 104 105
use FILL  FILL_254
timestamp 1554483974
transform 1 0 1624 0 -1 1370
box -8 -3 16 105
use FILL  FILL_255
timestamp 1554483974
transform 1 0 1632 0 -1 1370
box -8 -3 16 105
use NAND2X1  NAND2X1_7
timestamp 1554483974
transform 1 0 1640 0 -1 1370
box -8 -3 32 105
use OAI21X1  OAI21X1_7
timestamp 1554483974
transform -1 0 1696 0 -1 1370
box -8 -3 34 105
use FILL  FILL_256
timestamp 1554483974
transform 1 0 1696 0 -1 1370
box -8 -3 16 105
use FILL  FILL_258
timestamp 1554483974
transform 1 0 1704 0 -1 1370
box -8 -3 16 105
use FILL  FILL_260
timestamp 1554483974
transform 1 0 1712 0 -1 1370
box -8 -3 16 105
use FILL  FILL_262
timestamp 1554483974
transform 1 0 1720 0 -1 1370
box -8 -3 16 105
use FILL  FILL_264
timestamp 1554483974
transform 1 0 1728 0 -1 1370
box -8 -3 16 105
use FILL  FILL_266
timestamp 1554483974
transform 1 0 1736 0 -1 1370
box -8 -3 16 105
use FILL  FILL_268
timestamp 1554483974
transform 1 0 1744 0 -1 1370
box -8 -3 16 105
use FILL  FILL_270
timestamp 1554483974
transform 1 0 1752 0 -1 1370
box -8 -3 16 105
use FILL  FILL_272
timestamp 1554483974
transform 1 0 1760 0 -1 1370
box -8 -3 16 105
use FILL  FILL_274
timestamp 1554483974
transform 1 0 1768 0 -1 1370
box -8 -3 16 105
use UART_VIA1  UART_VIA1_7
timestamp 1554483974
transform 1 0 1825 0 1 1270
box -10 -3 10 3
use M2_M1  M2_M1_225
timestamp 1554483974
transform 1 0 196 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_235
timestamp 1554483974
transform 1 0 76 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_236
timestamp 1554483974
transform 1 0 132 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_237
timestamp 1554483974
transform 1 0 172 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_238
timestamp 1554483974
transform 1 0 180 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_239
timestamp 1554483974
transform 1 0 196 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_276
timestamp 1554483974
transform 1 0 156 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_277
timestamp 1554483974
transform 1 0 172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_243
timestamp 1554483974
transform 1 0 132 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_278
timestamp 1554483974
transform 1 0 196 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_279
timestamp 1554483974
transform 1 0 204 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_244
timestamp 1554483974
transform 1 0 196 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_280
timestamp 1554483974
transform 1 0 220 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_281
timestamp 1554483974
transform 1 0 236 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_317
timestamp 1554483974
transform 1 0 228 0 1 1195
box -2 -2 2 2
use M3_M2  M3_M2_225
timestamp 1554483974
transform 1 0 252 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_240
timestamp 1554483974
transform 1 0 252 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_282
timestamp 1554483974
transform 1 0 252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_241
timestamp 1554483974
transform 1 0 268 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_226
timestamp 1554483974
transform 1 0 284 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_254
timestamp 1554483974
transform 1 0 300 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_242
timestamp 1554483974
transform 1 0 324 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_243
timestamp 1554483974
transform 1 0 332 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_244
timestamp 1554483974
transform 1 0 348 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_245
timestamp 1554483974
transform 1 0 316 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_283
timestamp 1554483974
transform 1 0 332 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_284
timestamp 1554483974
transform 1 0 340 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_246
timestamp 1554483974
transform 1 0 332 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_255
timestamp 1554483974
transform 1 0 340 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_226
timestamp 1554483974
transform 1 0 436 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_245
timestamp 1554483974
transform 1 0 412 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_246
timestamp 1554483974
transform 1 0 420 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_247
timestamp 1554483974
transform 1 0 436 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_238
timestamp 1554483974
transform 1 0 452 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_248
timestamp 1554483974
transform 1 0 460 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_285
timestamp 1554483974
transform 1 0 444 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_286
timestamp 1554483974
transform 1 0 452 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_287
timestamp 1554483974
transform 1 0 468 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_288
timestamp 1554483974
transform 1 0 476 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_256
timestamp 1554483974
transform 1 0 412 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_247
timestamp 1554483974
transform 1 0 468 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_227
timestamp 1554483974
transform 1 0 516 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_249
timestamp 1554483974
transform 1 0 516 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_210
timestamp 1554483974
transform 1 0 556 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_214
timestamp 1554483974
transform 1 0 532 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_227
timestamp 1554483974
transform 1 0 532 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_289
timestamp 1554483974
transform 1 0 540 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_228
timestamp 1554483974
transform 1 0 564 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_250
timestamp 1554483974
transform 1 0 564 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_211
timestamp 1554483974
transform 1 0 596 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_215
timestamp 1554483974
transform 1 0 588 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_229
timestamp 1554483974
transform 1 0 588 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_290
timestamp 1554483974
transform 1 0 564 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_291
timestamp 1554483974
transform 1 0 572 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_248
timestamp 1554483974
transform 1 0 564 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_257
timestamp 1554483974
transform 1 0 556 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_216
timestamp 1554483974
transform 1 0 612 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_251
timestamp 1554483974
transform 1 0 612 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_228
timestamp 1554483974
transform 1 0 636 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_239
timestamp 1554483974
transform 1 0 628 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_252
timestamp 1554483974
transform 1 0 636 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_258
timestamp 1554483974
transform 1 0 620 0 1 1185
box -3 -3 3 3
use M2_M1  M2_M1_292
timestamp 1554483974
transform 1 0 636 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_249
timestamp 1554483974
transform 1 0 636 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_229
timestamp 1554483974
transform 1 0 692 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_253
timestamp 1554483974
transform 1 0 692 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_254
timestamp 1554483974
transform 1 0 708 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_293
timestamp 1554483974
transform 1 0 692 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_294
timestamp 1554483974
transform 1 0 700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_295
timestamp 1554483974
transform 1 0 716 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_259
timestamp 1554483974
transform 1 0 700 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_260
timestamp 1554483974
transform 1 0 724 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_250
timestamp 1554483974
transform 1 0 740 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_255
timestamp 1554483974
transform 1 0 772 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_296
timestamp 1554483974
transform 1 0 788 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_230
timestamp 1554483974
transform 1 0 812 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_256
timestamp 1554483974
transform 1 0 804 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_257
timestamp 1554483974
transform 1 0 820 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_297
timestamp 1554483974
transform 1 0 812 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_251
timestamp 1554483974
transform 1 0 804 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_217
timestamp 1554483974
transform 1 0 836 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_218
timestamp 1554483974
transform 1 0 892 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_258
timestamp 1554483974
transform 1 0 884 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_259
timestamp 1554483974
transform 1 0 892 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_298
timestamp 1554483974
transform 1 0 860 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_299
timestamp 1554483974
transform 1 0 916 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_300
timestamp 1554483974
transform 1 0 932 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_261
timestamp 1554483974
transform 1 0 940 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_252
timestamp 1554483974
transform 1 0 956 0 1 1195
box -3 -3 3 3
use M2_M1  M2_M1_230
timestamp 1554483974
transform 1 0 980 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_301
timestamp 1554483974
transform 1 0 996 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_253
timestamp 1554483974
transform 1 0 988 0 1 1195
box -3 -3 3 3
use M3_M2  M3_M2_231
timestamp 1554483974
transform 1 0 1012 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_232
timestamp 1554483974
transform 1 0 1060 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_260
timestamp 1554483974
transform 1 0 1036 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_240
timestamp 1554483974
transform 1 0 1044 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_302
timestamp 1554483974
transform 1 0 1012 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_261
timestamp 1554483974
transform 1 0 1100 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_303
timestamp 1554483974
transform 1 0 1060 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_304
timestamp 1554483974
transform 1 0 1068 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_262
timestamp 1554483974
transform 1 0 1020 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_263
timestamp 1554483974
transform 1 0 1044 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_233
timestamp 1554483974
transform 1 0 1124 0 1 1225
box -3 -3 3 3
use M3_M2  M3_M2_219
timestamp 1554483974
transform 1 0 1180 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_231
timestamp 1554483974
transform 1 0 1188 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_262
timestamp 1554483974
transform 1 0 1180 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_305
timestamp 1554483974
transform 1 0 1164 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_306
timestamp 1554483974
transform 1 0 1172 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_264
timestamp 1554483974
transform 1 0 1164 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_234
timestamp 1554483974
transform 1 0 1196 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_263
timestamp 1554483974
transform 1 0 1196 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_212
timestamp 1554483974
transform 1 0 1244 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_220
timestamp 1554483974
transform 1 0 1252 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_232
timestamp 1554483974
transform 1 0 1244 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_241
timestamp 1554483974
transform 1 0 1252 0 1 1215
box -3 -3 3 3
use M2_M1  M2_M1_307
timestamp 1554483974
transform 1 0 1252 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_264
timestamp 1554483974
transform 1 0 1268 0 1 1215
box -2 -2 2 2
use M3_M2  M3_M2_265
timestamp 1554483974
transform 1 0 1268 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_208
timestamp 1554483974
transform 1 0 1348 0 1 1255
box -3 -3 3 3
use M3_M2  M3_M2_213
timestamp 1554483974
transform 1 0 1340 0 1 1245
box -3 -3 3 3
use M3_M2  M3_M2_221
timestamp 1554483974
transform 1 0 1316 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_233
timestamp 1554483974
transform 1 0 1316 0 1 1225
box -2 -2 2 2
use M3_M2  M3_M2_242
timestamp 1554483974
transform 1 0 1324 0 1 1215
box -3 -3 3 3
use M3_M2  M3_M2_222
timestamp 1554483974
transform 1 0 1372 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_235
timestamp 1554483974
transform 1 0 1396 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_265
timestamp 1554483974
transform 1 0 1340 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_266
timestamp 1554483974
transform 1 0 1356 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_267
timestamp 1554483974
transform 1 0 1372 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_268
timestamp 1554483974
transform 1 0 1388 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_308
timestamp 1554483974
transform 1 0 1324 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_309
timestamp 1554483974
transform 1 0 1364 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_209
timestamp 1554483974
transform 1 0 1420 0 1 1255
box -3 -3 3 3
use M2_M1  M2_M1_310
timestamp 1554483974
transform 1 0 1412 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_266
timestamp 1554483974
transform 1 0 1412 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_236
timestamp 1554483974
transform 1 0 1508 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_269
timestamp 1554483974
transform 1 0 1476 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_270
timestamp 1554483974
transform 1 0 1508 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_271
timestamp 1554483974
transform 1 0 1516 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_272
timestamp 1554483974
transform 1 0 1524 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_273
timestamp 1554483974
transform 1 0 1532 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_311
timestamp 1554483974
transform 1 0 1428 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_312
timestamp 1554483974
transform 1 0 1516 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_267
timestamp 1554483974
transform 1 0 1532 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_223
timestamp 1554483974
transform 1 0 1604 0 1 1235
box -3 -3 3 3
use M2_M1  M2_M1_274
timestamp 1554483974
transform 1 0 1604 0 1 1215
box -2 -2 2 2
use M2_M1  M2_M1_313
timestamp 1554483974
transform 1 0 1628 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_314
timestamp 1554483974
transform 1 0 1644 0 1 1205
box -2 -2 2 2
use M3_M2  M3_M2_268
timestamp 1554483974
transform 1 0 1644 0 1 1185
box -3 -3 3 3
use M3_M2  M3_M2_224
timestamp 1554483974
transform 1 0 1676 0 1 1235
box -3 -3 3 3
use M3_M2  M3_M2_237
timestamp 1554483974
transform 1 0 1660 0 1 1225
box -3 -3 3 3
use M2_M1  M2_M1_234
timestamp 1554483974
transform 1 0 1668 0 1 1225
box -2 -2 2 2
use M2_M1  M2_M1_315
timestamp 1554483974
transform 1 0 1676 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_316
timestamp 1554483974
transform 1 0 1700 0 1 1205
box -2 -2 2 2
use M2_M1  M2_M1_275
timestamp 1554483974
transform 1 0 1732 0 1 1215
box -2 -2 2 2
use UART_VIA1  UART_VIA1_8
timestamp 1554483974
transform 1 0 48 0 1 1170
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_8
timestamp 1554483974
transform -1 0 168 0 1 1170
box -8 -3 104 105
use OAI21X1  OAI21X1_8
timestamp 1554483974
transform 1 0 168 0 1 1170
box -8 -3 34 105
use INVX2  INVX2_10
timestamp 1554483974
transform 1 0 200 0 1 1170
box -9 -3 26 105
use FILL  FILL_275
timestamp 1554483974
transform 1 0 216 0 1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_5
timestamp 1554483974
transform 1 0 224 0 1 1170
box -8 -3 32 105
use FILL  FILL_276
timestamp 1554483974
transform 1 0 248 0 1 1170
box -8 -3 16 105
use FILL  FILL_291
timestamp 1554483974
transform 1 0 256 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_8
timestamp 1554483974
transform 1 0 264 0 1 1170
box -8 -3 32 105
use FILL  FILL_293
timestamp 1554483974
transform 1 0 288 0 1 1170
box -8 -3 16 105
use FILL  FILL_298
timestamp 1554483974
transform 1 0 296 0 1 1170
box -8 -3 16 105
use FILL  FILL_300
timestamp 1554483974
transform 1 0 304 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_269
timestamp 1554483974
transform 1 0 340 0 1 1175
box -3 -3 3 3
use NAND2X1  NAND2X1_9
timestamp 1554483974
transform -1 0 336 0 1 1170
box -8 -3 32 105
use INVX2  INVX2_12
timestamp 1554483974
transform 1 0 336 0 1 1170
box -9 -3 26 105
use FILL  FILL_301
timestamp 1554483974
transform 1 0 352 0 1 1170
box -8 -3 16 105
use FILL  FILL_305
timestamp 1554483974
transform 1 0 360 0 1 1170
box -8 -3 16 105
use FILL  FILL_307
timestamp 1554483974
transform 1 0 368 0 1 1170
box -8 -3 16 105
use FILL  FILL_309
timestamp 1554483974
transform 1 0 376 0 1 1170
box -8 -3 16 105
use FILL  FILL_311
timestamp 1554483974
transform 1 0 384 0 1 1170
box -8 -3 16 105
use FILL  FILL_313
timestamp 1554483974
transform 1 0 392 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_270
timestamp 1554483974
transform 1 0 420 0 1 1175
box -3 -3 3 3
use NAND2X1  NAND2X1_10
timestamp 1554483974
transform 1 0 400 0 1 1170
box -8 -3 32 105
use INVX2  INVX2_13
timestamp 1554483974
transform -1 0 440 0 1 1170
box -9 -3 26 105
use AOI22X1  AOI22X1_3
timestamp 1554483974
transform 1 0 440 0 1 1170
box -8 -3 46 105
use FILL  FILL_315
timestamp 1554483974
transform 1 0 480 0 1 1170
box -8 -3 16 105
use FILL  FILL_316
timestamp 1554483974
transform 1 0 488 0 1 1170
box -8 -3 16 105
use FILL  FILL_317
timestamp 1554483974
transform 1 0 496 0 1 1170
box -8 -3 16 105
use FILL  FILL_319
timestamp 1554483974
transform 1 0 504 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_11
timestamp 1554483974
transform 1 0 512 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_10
timestamp 1554483974
transform 1 0 536 0 1 1170
box -8 -3 34 105
use NAND2X1  NAND2X1_12
timestamp 1554483974
transform 1 0 568 0 1 1170
box -8 -3 32 105
use FILL  FILL_324
timestamp 1554483974
transform 1 0 592 0 1 1170
box -8 -3 16 105
use FILL  FILL_329
timestamp 1554483974
transform 1 0 600 0 1 1170
box -8 -3 16 105
use FILL  FILL_330
timestamp 1554483974
transform 1 0 608 0 1 1170
box -8 -3 16 105
use FILL  FILL_331
timestamp 1554483974
transform 1 0 616 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_14
timestamp 1554483974
transform -1 0 640 0 1 1170
box -9 -3 26 105
use FILL  FILL_332
timestamp 1554483974
transform 1 0 640 0 1 1170
box -8 -3 16 105
use INVX2  INVX2_15
timestamp 1554483974
transform -1 0 664 0 1 1170
box -9 -3 26 105
use FILL  FILL_333
timestamp 1554483974
transform 1 0 664 0 1 1170
box -8 -3 16 105
use FILL  FILL_334
timestamp 1554483974
transform 1 0 672 0 1 1170
box -8 -3 16 105
use FILL  FILL_335
timestamp 1554483974
transform 1 0 680 0 1 1170
box -8 -3 16 105
use AOI22X1  AOI22X1_4
timestamp 1554483974
transform -1 0 728 0 1 1170
box -8 -3 46 105
use FILL  FILL_336
timestamp 1554483974
transform 1 0 728 0 1 1170
box -8 -3 16 105
use FILL  FILL_337
timestamp 1554483974
transform 1 0 736 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_271
timestamp 1554483974
transform 1 0 756 0 1 1175
box -3 -3 3 3
use FILL  FILL_338
timestamp 1554483974
transform 1 0 744 0 1 1170
box -8 -3 16 105
use FILL  FILL_339
timestamp 1554483974
transform 1 0 752 0 1 1170
box -8 -3 16 105
use FILL  FILL_340
timestamp 1554483974
transform 1 0 760 0 1 1170
box -8 -3 16 105
use FILL  FILL_341
timestamp 1554483974
transform 1 0 768 0 1 1170
box -8 -3 16 105
use FILL  FILL_342
timestamp 1554483974
transform 1 0 776 0 1 1170
box -8 -3 16 105
use FILL  FILL_343
timestamp 1554483974
transform 1 0 784 0 1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_4
timestamp 1554483974
transform -1 0 832 0 1 1170
box -8 -3 46 105
use FILL  FILL_344
timestamp 1554483974
transform 1 0 832 0 1 1170
box -8 -3 16 105
use FILL  FILL_345
timestamp 1554483974
transform 1 0 840 0 1 1170
box -8 -3 16 105
use FILL  FILL_346
timestamp 1554483974
transform 1 0 848 0 1 1170
box -8 -3 16 105
use XOR2X1  XOR2X1_5
timestamp 1554483974
transform 1 0 856 0 1 1170
box -8 -3 64 105
use FILL  FILL_347
timestamp 1554483974
transform 1 0 912 0 1 1170
box -8 -3 16 105
use FILL  FILL_351
timestamp 1554483974
transform 1 0 920 0 1 1170
box -8 -3 16 105
use FILL  FILL_353
timestamp 1554483974
transform 1 0 928 0 1 1170
box -8 -3 16 105
use FILL  FILL_354
timestamp 1554483974
transform 1 0 936 0 1 1170
box -8 -3 16 105
use FILL  FILL_355
timestamp 1554483974
transform 1 0 944 0 1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_13
timestamp 1554483974
transform 1 0 952 0 1 1170
box -8 -3 34 105
use FILL  FILL_356
timestamp 1554483974
transform 1 0 984 0 1 1170
box -8 -3 16 105
use FILL  FILL_357
timestamp 1554483974
transform 1 0 992 0 1 1170
box -8 -3 16 105
use FILL  FILL_358
timestamp 1554483974
transform 1 0 1000 0 1 1170
box -8 -3 16 105
use M3_M2  M3_M2_272
timestamp 1554483974
transform 1 0 1068 0 1 1175
box -3 -3 3 3
use XOR2X1  XOR2X1_8
timestamp 1554483974
transform 1 0 1008 0 1 1170
box -8 -3 64 105
use XNOR2X1  XNOR2X1_3
timestamp 1554483974
transform 1 0 1064 0 1 1170
box -8 -3 64 105
use FILL  FILL_359
timestamp 1554483974
transform 1 0 1120 0 1 1170
box -8 -3 16 105
use FILL  FILL_360
timestamp 1554483974
transform 1 0 1128 0 1 1170
box -8 -3 16 105
use FILL  FILL_361
timestamp 1554483974
transform 1 0 1136 0 1 1170
box -8 -3 16 105
use FILL  FILL_362
timestamp 1554483974
transform 1 0 1144 0 1 1170
box -8 -3 16 105
use FILL  FILL_363
timestamp 1554483974
transform 1 0 1152 0 1 1170
box -8 -3 16 105
use FILL  FILL_366
timestamp 1554483974
transform 1 0 1160 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_14
timestamp 1554483974
transform 1 0 1168 0 1 1170
box -8 -3 32 105
use FILL  FILL_368
timestamp 1554483974
transform 1 0 1192 0 1 1170
box -8 -3 16 105
use FILL  FILL_369
timestamp 1554483974
transform 1 0 1200 0 1 1170
box -8 -3 16 105
use LATCH  LATCH_6
timestamp 1554483974
transform -1 0 1264 0 1 1170
box -8 -3 64 105
use FILL  FILL_370
timestamp 1554483974
transform 1 0 1264 0 1 1170
box -8 -3 16 105
use FILL  FILL_371
timestamp 1554483974
transform 1 0 1272 0 1 1170
box -8 -3 16 105
use LATCH  LATCH_7
timestamp 1554483974
transform -1 0 1336 0 1 1170
box -8 -3 64 105
use AND2X2  AND2X2_6
timestamp 1554483974
transform -1 0 1368 0 1 1170
box -8 -3 40 105
use AND2X2  AND2X2_7
timestamp 1554483974
transform -1 0 1400 0 1 1170
box -8 -3 40 105
use FILL  FILL_372
timestamp 1554483974
transform 1 0 1400 0 1 1170
box -8 -3 16 105
use FILL  FILL_382
timestamp 1554483974
transform 1 0 1408 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_14
timestamp 1554483974
transform 1 0 1416 0 1 1170
box -8 -3 104 105
use INVX2  INVX2_17
timestamp 1554483974
transform 1 0 1512 0 1 1170
box -9 -3 26 105
use FILL  FILL_384
timestamp 1554483974
transform 1 0 1528 0 1 1170
box -8 -3 16 105
use FILL  FILL_391
timestamp 1554483974
transform 1 0 1536 0 1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_15
timestamp 1554483974
transform -1 0 1640 0 1 1170
box -8 -3 104 105
use FILL  FILL_392
timestamp 1554483974
transform 1 0 1640 0 1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_18
timestamp 1554483974
transform 1 0 1648 0 1 1170
box -8 -3 32 105
use OAI21X1  OAI21X1_14
timestamp 1554483974
transform -1 0 1704 0 1 1170
box -8 -3 34 105
use FILL  FILL_393
timestamp 1554483974
transform 1 0 1704 0 1 1170
box -8 -3 16 105
use FILL  FILL_394
timestamp 1554483974
transform 1 0 1712 0 1 1170
box -8 -3 16 105
use FILL  FILL_395
timestamp 1554483974
transform 1 0 1720 0 1 1170
box -8 -3 16 105
use FILL  FILL_401
timestamp 1554483974
transform 1 0 1728 0 1 1170
box -8 -3 16 105
use FILL  FILL_403
timestamp 1554483974
transform 1 0 1736 0 1 1170
box -8 -3 16 105
use FILL  FILL_404
timestamp 1554483974
transform 1 0 1744 0 1 1170
box -8 -3 16 105
use FILL  FILL_405
timestamp 1554483974
transform 1 0 1752 0 1 1170
box -8 -3 16 105
use FILL  FILL_407
timestamp 1554483974
transform 1 0 1760 0 1 1170
box -8 -3 16 105
use FILL  FILL_409
timestamp 1554483974
transform 1 0 1768 0 1 1170
box -8 -3 16 105
use UART_VIA1  UART_VIA1_9
timestamp 1554483974
transform 1 0 1801 0 1 1170
box -10 -3 10 3
use M3_M2  M3_M2_286
timestamp 1554483974
transform 1 0 76 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_318
timestamp 1554483974
transform 1 0 100 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_287
timestamp 1554483974
transform 1 0 108 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_321
timestamp 1554483974
transform 1 0 124 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_288
timestamp 1554483974
transform 1 0 140 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_322
timestamp 1554483974
transform 1 0 156 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_353
timestamp 1554483974
transform 1 0 156 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_316
timestamp 1554483974
transform 1 0 156 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_323
timestamp 1554483974
transform 1 0 172 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_354
timestamp 1554483974
transform 1 0 180 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_289
timestamp 1554483974
transform 1 0 204 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_300
timestamp 1554483974
transform 1 0 212 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_355
timestamp 1554483974
transform 1 0 236 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_356
timestamp 1554483974
transform 1 0 244 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_387
timestamp 1554483974
transform 1 0 220 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_317
timestamp 1554483974
transform 1 0 236 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_324
timestamp 1554483974
transform 1 0 220 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_275
timestamp 1554483974
transform 1 0 284 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_319
timestamp 1554483974
transform 1 0 284 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_301
timestamp 1554483974
transform 1 0 284 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_324
timestamp 1554483974
transform 1 0 300 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_357
timestamp 1554483974
transform 1 0 292 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_325
timestamp 1554483974
transform 1 0 292 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_318
timestamp 1554483974
transform 1 0 308 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_325
timestamp 1554483974
transform 1 0 348 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_358
timestamp 1554483974
transform 1 0 348 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_331
timestamp 1554483974
transform 1 0 348 0 1 1095
box -3 -3 3 3
use M3_M2  M3_M2_276
timestamp 1554483974
transform 1 0 492 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_326
timestamp 1554483974
transform 1 0 412 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_359
timestamp 1554483974
transform 1 0 436 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_360
timestamp 1554483974
transform 1 0 492 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_319
timestamp 1554483974
transform 1 0 436 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_332
timestamp 1554483974
transform 1 0 476 0 1 1095
box -3 -3 3 3
use M2_M1  M2_M1_327
timestamp 1554483974
transform 1 0 540 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_361
timestamp 1554483974
transform 1 0 548 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_277
timestamp 1554483974
transform 1 0 572 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_328
timestamp 1554483974
transform 1 0 572 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_388
timestamp 1554483974
transform 1 0 580 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_290
timestamp 1554483974
transform 1 0 644 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_329
timestamp 1554483974
transform 1 0 612 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_330
timestamp 1554483974
transform 1 0 628 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_331
timestamp 1554483974
transform 1 0 644 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_332
timestamp 1554483974
transform 1 0 652 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_310
timestamp 1554483974
transform 1 0 604 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_389
timestamp 1554483974
transform 1 0 596 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_362
timestamp 1554483974
transform 1 0 620 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_363
timestamp 1554483974
transform 1 0 636 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_311
timestamp 1554483974
transform 1 0 652 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_291
timestamp 1554483974
transform 1 0 708 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_333
timestamp 1554483974
transform 1 0 700 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_334
timestamp 1554483974
transform 1 0 708 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_278
timestamp 1554483974
transform 1 0 772 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_279
timestamp 1554483974
transform 1 0 828 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_292
timestamp 1554483974
transform 1 0 764 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_293
timestamp 1554483974
transform 1 0 860 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_335
timestamp 1554483974
transform 1 0 756 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_336
timestamp 1554483974
transform 1 0 844 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_337
timestamp 1554483974
transform 1 0 860 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_364
timestamp 1554483974
transform 1 0 700 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_365
timestamp 1554483974
transform 1 0 732 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_366
timestamp 1554483974
transform 1 0 764 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_367
timestamp 1554483974
transform 1 0 812 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_312
timestamp 1554483974
transform 1 0 820 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_326
timestamp 1554483974
transform 1 0 844 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_302
timestamp 1554483974
transform 1 0 868 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_338
timestamp 1554483974
transform 1 0 876 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_303
timestamp 1554483974
transform 1 0 892 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_368
timestamp 1554483974
transform 1 0 868 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_313
timestamp 1554483974
transform 1 0 876 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_369
timestamp 1554483974
transform 1 0 892 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_390
timestamp 1554483974
transform 1 0 876 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_391
timestamp 1554483974
transform 1 0 916 0 1 1115
box -2 -2 2 2
use M2_M1  M2_M1_339
timestamp 1554483974
transform 1 0 932 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_304
timestamp 1554483974
transform 1 0 948 0 1 1135
box -3 -3 3 3
use M3_M2  M3_M2_294
timestamp 1554483974
transform 1 0 1044 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_340
timestamp 1554483974
transform 1 0 956 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_305
timestamp 1554483974
transform 1 0 980 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_341
timestamp 1554483974
transform 1 0 1044 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_370
timestamp 1554483974
transform 1 0 948 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_371
timestamp 1554483974
transform 1 0 956 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_372
timestamp 1554483974
transform 1 0 996 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_280
timestamp 1554483974
transform 1 0 1068 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_295
timestamp 1554483974
transform 1 0 1068 0 1 1145
box -3 -3 3 3
use M3_M2  M3_M2_296
timestamp 1554483974
transform 1 0 1148 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_342
timestamp 1554483974
transform 1 0 1068 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_373
timestamp 1554483974
transform 1 0 1116 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_327
timestamp 1554483974
transform 1 0 1100 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_374
timestamp 1554483974
transform 1 0 1156 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_297
timestamp 1554483974
transform 1 0 1172 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_375
timestamp 1554483974
transform 1 0 1196 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_392
timestamp 1554483974
transform 1 0 1204 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_328
timestamp 1554483974
transform 1 0 1204 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_343
timestamp 1554483974
transform 1 0 1220 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_376
timestamp 1554483974
transform 1 0 1236 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_281
timestamp 1554483974
transform 1 0 1268 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_344
timestamp 1554483974
transform 1 0 1268 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_345
timestamp 1554483974
transform 1 0 1356 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_377
timestamp 1554483974
transform 1 0 1316 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_378
timestamp 1554483974
transform 1 0 1364 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_393
timestamp 1554483974
transform 1 0 1252 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_320
timestamp 1554483974
transform 1 0 1316 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_321
timestamp 1554483974
transform 1 0 1356 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_329
timestamp 1554483974
transform 1 0 1252 0 1 1105
box -3 -3 3 3
use M3_M2  M3_M2_282
timestamp 1554483974
transform 1 0 1380 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_394
timestamp 1554483974
transform 1 0 1372 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_330
timestamp 1554483974
transform 1 0 1372 0 1 1105
box -3 -3 3 3
use M2_M1  M2_M1_379
timestamp 1554483974
transform 1 0 1404 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_395
timestamp 1554483974
transform 1 0 1396 0 1 1115
box -2 -2 2 2
use M3_M2  M3_M2_283
timestamp 1554483974
transform 1 0 1428 0 1 1155
box -3 -3 3 3
use M2_M1  M2_M1_320
timestamp 1554483974
transform 1 0 1444 0 1 1145
box -2 -2 2 2
use M3_M2  M3_M2_322
timestamp 1554483974
transform 1 0 1444 0 1 1115
box -3 -3 3 3
use M2_M1  M2_M1_346
timestamp 1554483974
transform 1 0 1460 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_273
timestamp 1554483974
transform 1 0 1476 0 1 1165
box -3 -3 3 3
use M3_M2  M3_M2_306
timestamp 1554483974
transform 1 0 1468 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_380
timestamp 1554483974
transform 1 0 1476 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_274
timestamp 1554483974
transform 1 0 1508 0 1 1165
box -3 -3 3 3
use M2_M1  M2_M1_347
timestamp 1554483974
transform 1 0 1508 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_307
timestamp 1554483974
transform 1 0 1516 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_348
timestamp 1554483974
transform 1 0 1524 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_381
timestamp 1554483974
transform 1 0 1500 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_382
timestamp 1554483974
transform 1 0 1516 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_323
timestamp 1554483974
transform 1 0 1516 0 1 1115
box -3 -3 3 3
use M3_M2  M3_M2_284
timestamp 1554483974
transform 1 0 1580 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_285
timestamp 1554483974
transform 1 0 1628 0 1 1155
box -3 -3 3 3
use M3_M2  M3_M2_298
timestamp 1554483974
transform 1 0 1628 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_349
timestamp 1554483974
transform 1 0 1580 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_383
timestamp 1554483974
transform 1 0 1628 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_299
timestamp 1554483974
transform 1 0 1700 0 1 1145
box -3 -3 3 3
use M2_M1  M2_M1_350
timestamp 1554483974
transform 1 0 1684 0 1 1135
box -2 -2 2 2
use M2_M1  M2_M1_351
timestamp 1554483974
transform 1 0 1700 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_308
timestamp 1554483974
transform 1 0 1708 0 1 1135
box -3 -3 3 3
use M2_M1  M2_M1_384
timestamp 1554483974
transform 1 0 1676 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_385
timestamp 1554483974
transform 1 0 1692 0 1 1125
box -2 -2 2 2
use M3_M2  M3_M2_314
timestamp 1554483974
transform 1 0 1700 0 1 1125
box -3 -3 3 3
use M2_M1  M2_M1_386
timestamp 1554483974
transform 1 0 1708 0 1 1125
box -2 -2 2 2
use M2_M1  M2_M1_352
timestamp 1554483974
transform 1 0 1724 0 1 1135
box -2 -2 2 2
use M3_M2  M3_M2_315
timestamp 1554483974
transform 1 0 1724 0 1 1125
box -3 -3 3 3
use M3_M2  M3_M2_309
timestamp 1554483974
transform 1 0 1740 0 1 1135
box -3 -3 3 3
use UART_VIA1  UART_VIA1_10
timestamp 1554483974
transform 1 0 24 0 1 1070
box -10 -3 10 3
use FILL  FILL_277
timestamp 1554483974
transform 1 0 72 0 -1 1170
box -8 -3 16 105
use FILL  FILL_278
timestamp 1554483974
transform 1 0 80 0 -1 1170
box -8 -3 16 105
use FILL  FILL_279
timestamp 1554483974
transform 1 0 88 0 -1 1170
box -8 -3 16 105
use NOR2X1  NOR2X1_6
timestamp 1554483974
transform 1 0 96 0 -1 1170
box -8 -3 32 105
use FILL  FILL_280
timestamp 1554483974
transform 1 0 120 0 -1 1170
box -8 -3 16 105
use FILL  FILL_281
timestamp 1554483974
transform 1 0 128 0 -1 1170
box -8 -3 16 105
use FILL  FILL_282
timestamp 1554483974
transform 1 0 136 0 -1 1170
box -8 -3 16 105
use FILL  FILL_283
timestamp 1554483974
transform 1 0 144 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_11
timestamp 1554483974
transform 1 0 152 0 -1 1170
box -9 -3 26 105
use FILL  FILL_284
timestamp 1554483974
transform 1 0 168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_285
timestamp 1554483974
transform 1 0 176 0 -1 1170
box -8 -3 16 105
use FILL  FILL_286
timestamp 1554483974
transform 1 0 184 0 -1 1170
box -8 -3 16 105
use FILL  FILL_287
timestamp 1554483974
transform 1 0 192 0 -1 1170
box -8 -3 16 105
use FILL  FILL_288
timestamp 1554483974
transform 1 0 200 0 -1 1170
box -8 -3 16 105
use FILL  FILL_289
timestamp 1554483974
transform 1 0 208 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_9
timestamp 1554483974
transform -1 0 248 0 -1 1170
box -8 -3 34 105
use FILL  FILL_290
timestamp 1554483974
transform 1 0 248 0 -1 1170
box -8 -3 16 105
use FILL  FILL_292
timestamp 1554483974
transform 1 0 256 0 -1 1170
box -8 -3 16 105
use FILL  FILL_294
timestamp 1554483974
transform 1 0 264 0 -1 1170
box -8 -3 16 105
use FILL  FILL_295
timestamp 1554483974
transform 1 0 272 0 -1 1170
box -8 -3 16 105
use FILL  FILL_296
timestamp 1554483974
transform 1 0 280 0 -1 1170
box -8 -3 16 105
use FILL  FILL_297
timestamp 1554483974
transform 1 0 288 0 -1 1170
box -8 -3 16 105
use FILL  FILL_299
timestamp 1554483974
transform 1 0 296 0 -1 1170
box -8 -3 16 105
use FILL  FILL_302
timestamp 1554483974
transform 1 0 304 0 -1 1170
box -8 -3 16 105
use FILL  FILL_303
timestamp 1554483974
transform 1 0 312 0 -1 1170
box -8 -3 16 105
use AOI21X1  AOI21X1_0
timestamp 1554483974
transform -1 0 352 0 -1 1170
box -7 -3 39 105
use FILL  FILL_304
timestamp 1554483974
transform 1 0 352 0 -1 1170
box -8 -3 16 105
use FILL  FILL_306
timestamp 1554483974
transform 1 0 360 0 -1 1170
box -8 -3 16 105
use FILL  FILL_308
timestamp 1554483974
transform 1 0 368 0 -1 1170
box -8 -3 16 105
use FILL  FILL_310
timestamp 1554483974
transform 1 0 376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_312
timestamp 1554483974
transform 1 0 384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_314
timestamp 1554483974
transform 1 0 392 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_9
timestamp 1554483974
transform 1 0 400 0 -1 1170
box -8 -3 104 105
use FILL  FILL_318
timestamp 1554483974
transform 1 0 496 0 -1 1170
box -8 -3 16 105
use FILL  FILL_320
timestamp 1554483974
transform 1 0 504 0 -1 1170
box -8 -3 16 105
use FILL  FILL_321
timestamp 1554483974
transform 1 0 512 0 -1 1170
box -8 -3 16 105
use FILL  FILL_322
timestamp 1554483974
transform 1 0 520 0 -1 1170
box -8 -3 16 105
use FILL  FILL_323
timestamp 1554483974
transform 1 0 528 0 -1 1170
box -8 -3 16 105
use OAI21X1  OAI21X1_11
timestamp 1554483974
transform 1 0 536 0 -1 1170
box -8 -3 34 105
use FILL  FILL_325
timestamp 1554483974
transform 1 0 568 0 -1 1170
box -8 -3 16 105
use FILL  FILL_326
timestamp 1554483974
transform 1 0 576 0 -1 1170
box -8 -3 16 105
use FILL  FILL_327
timestamp 1554483974
transform 1 0 584 0 -1 1170
box -8 -3 16 105
use FILL  FILL_328
timestamp 1554483974
transform 1 0 592 0 -1 1170
box -8 -3 16 105
use FILL  FILL_348
timestamp 1554483974
transform 1 0 600 0 -1 1170
box -8 -3 16 105
use OAI22X1  OAI22X1_5
timestamp 1554483974
transform -1 0 648 0 -1 1170
box -8 -3 46 105
use XOR2X1  XOR2X1_6
timestamp 1554483974
transform 1 0 648 0 -1 1170
box -8 -3 64 105
use XOR2X1  XOR2X1_7
timestamp 1554483974
transform 1 0 704 0 -1 1170
box -8 -3 64 105
use DFFNEGX1  DFFNEGX1_10
timestamp 1554483974
transform -1 0 856 0 -1 1170
box -8 -3 104 105
use INVX2  INVX2_16
timestamp 1554483974
transform 1 0 856 0 -1 1170
box -9 -3 26 105
use OAI21X1  OAI21X1_12
timestamp 1554483974
transform -1 0 904 0 -1 1170
box -8 -3 34 105
use FILL  FILL_349
timestamp 1554483974
transform 1 0 904 0 -1 1170
box -8 -3 16 105
use FILL  FILL_350
timestamp 1554483974
transform 1 0 912 0 -1 1170
box -8 -3 16 105
use FILL  FILL_352
timestamp 1554483974
transform 1 0 920 0 -1 1170
box -8 -3 16 105
use FILL  FILL_364
timestamp 1554483974
transform 1 0 928 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_13
timestamp 1554483974
transform -1 0 960 0 -1 1170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_11
timestamp 1554483974
transform -1 0 1056 0 -1 1170
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_12
timestamp 1554483974
transform 1 0 1056 0 -1 1170
box -8 -3 104 105
use FILL  FILL_365
timestamp 1554483974
transform 1 0 1152 0 -1 1170
box -8 -3 16 105
use FILL  FILL_367
timestamp 1554483974
transform 1 0 1160 0 -1 1170
box -8 -3 16 105
use FILL  FILL_373
timestamp 1554483974
transform 1 0 1168 0 -1 1170
box -8 -3 16 105
use FILL  FILL_374
timestamp 1554483974
transform 1 0 1176 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_15
timestamp 1554483974
transform 1 0 1184 0 -1 1170
box -8 -3 32 105
use FILL  FILL_375
timestamp 1554483974
transform 1 0 1208 0 -1 1170
box -8 -3 16 105
use FILL  FILL_376
timestamp 1554483974
transform 1 0 1216 0 -1 1170
box -8 -3 16 105
use FILL  FILL_377
timestamp 1554483974
transform 1 0 1224 0 -1 1170
box -8 -3 16 105
use NAND2X1  NAND2X1_16
timestamp 1554483974
transform 1 0 1232 0 -1 1170
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_13
timestamp 1554483974
transform 1 0 1256 0 -1 1170
box -8 -3 104 105
use NAND2X1  NAND2X1_17
timestamp 1554483974
transform 1 0 1352 0 -1 1170
box -8 -3 32 105
use FILL  FILL_378
timestamp 1554483974
transform 1 0 1376 0 -1 1170
box -8 -3 16 105
use FILL  FILL_379
timestamp 1554483974
transform 1 0 1384 0 -1 1170
box -8 -3 16 105
use FILL  FILL_380
timestamp 1554483974
transform 1 0 1392 0 -1 1170
box -8 -3 16 105
use FILL  FILL_381
timestamp 1554483974
transform 1 0 1400 0 -1 1170
box -8 -3 16 105
use FILL  FILL_383
timestamp 1554483974
transform 1 0 1408 0 -1 1170
box -8 -3 16 105
use FILL  FILL_385
timestamp 1554483974
transform 1 0 1416 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_18
timestamp 1554483974
transform -1 0 1440 0 -1 1170
box -9 -3 26 105
use FILL  FILL_386
timestamp 1554483974
transform 1 0 1440 0 -1 1170
box -8 -3 16 105
use FILL  FILL_387
timestamp 1554483974
transform 1 0 1448 0 -1 1170
box -8 -3 16 105
use FILL  FILL_388
timestamp 1554483974
transform 1 0 1456 0 -1 1170
box -8 -3 16 105
use FILL  FILL_389
timestamp 1554483974
transform 1 0 1464 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_19
timestamp 1554483974
transform 1 0 1472 0 -1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_6
timestamp 1554483974
transform 1 0 1488 0 -1 1170
box -8 -3 46 105
use FILL  FILL_390
timestamp 1554483974
transform 1 0 1528 0 -1 1170
box -8 -3 16 105
use FILL  FILL_396
timestamp 1554483974
transform 1 0 1536 0 -1 1170
box -8 -3 16 105
use FILL  FILL_397
timestamp 1554483974
transform 1 0 1544 0 -1 1170
box -8 -3 16 105
use M3_M2  M3_M2_333
timestamp 1554483974
transform 1 0 1564 0 1 1075
box -3 -3 3 3
use FILL  FILL_398
timestamp 1554483974
transform 1 0 1552 0 -1 1170
box -8 -3 16 105
use FILL  FILL_399
timestamp 1554483974
transform 1 0 1560 0 -1 1170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_16
timestamp 1554483974
transform 1 0 1568 0 -1 1170
box -8 -3 104 105
use M3_M2  M3_M2_334
timestamp 1554483974
transform 1 0 1676 0 1 1075
box -3 -3 3 3
use INVX2  INVX2_20
timestamp 1554483974
transform 1 0 1664 0 -1 1170
box -9 -3 26 105
use OAI22X1  OAI22X1_7
timestamp 1554483974
transform -1 0 1720 0 -1 1170
box -8 -3 46 105
use FILL  FILL_400
timestamp 1554483974
transform 1 0 1720 0 -1 1170
box -8 -3 16 105
use FILL  FILL_402
timestamp 1554483974
transform 1 0 1728 0 -1 1170
box -8 -3 16 105
use INVX2  INVX2_21
timestamp 1554483974
transform 1 0 1736 0 -1 1170
box -9 -3 26 105
use FILL  FILL_406
timestamp 1554483974
transform 1 0 1752 0 -1 1170
box -8 -3 16 105
use FILL  FILL_408
timestamp 1554483974
transform 1 0 1760 0 -1 1170
box -8 -3 16 105
use FILL  FILL_410
timestamp 1554483974
transform 1 0 1768 0 -1 1170
box -8 -3 16 105
use UART_VIA1  UART_VIA1_11
timestamp 1554483974
transform 1 0 1825 0 1 1070
box -10 -3 10 3
use M2_M1  M2_M1_396
timestamp 1554483974
transform 1 0 124 0 1 1035
box -2 -2 2 2
use M2_M1  M2_M1_397
timestamp 1554483974
transform 1 0 108 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_407
timestamp 1554483974
transform 1 0 124 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_445
timestamp 1554483974
transform 1 0 140 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_482
timestamp 1554483974
transform 1 0 140 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_335
timestamp 1554483974
transform 1 0 164 0 1 1055
box -3 -3 3 3
use M2_M1  M2_M1_398
timestamp 1554483974
transform 1 0 156 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_352
timestamp 1554483974
transform 1 0 156 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_361
timestamp 1554483974
transform 1 0 156 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_483
timestamp 1554483974
transform 1 0 164 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_339
timestamp 1554483974
transform 1 0 188 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_408
timestamp 1554483974
transform 1 0 188 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_353
timestamp 1554483974
transform 1 0 196 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_446
timestamp 1554483974
transform 1 0 196 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_409
timestamp 1554483974
transform 1 0 212 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_484
timestamp 1554483974
transform 1 0 228 0 1 995
box -2 -2 2 2
use M3_M2  M3_M2_354
timestamp 1554483974
transform 1 0 252 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_447
timestamp 1554483974
transform 1 0 276 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_410
timestamp 1554483974
transform 1 0 284 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_336
timestamp 1554483974
transform 1 0 324 0 1 1055
box -3 -3 3 3
use M3_M2  M3_M2_337
timestamp 1554483974
transform 1 0 324 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_338
timestamp 1554483974
transform 1 0 348 0 1 1045
box -3 -3 3 3
use M3_M2  M3_M2_340
timestamp 1554483974
transform 1 0 332 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_411
timestamp 1554483974
transform 1 0 300 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_412
timestamp 1554483974
transform 1 0 316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_413
timestamp 1554483974
transform 1 0 332 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_448
timestamp 1554483974
transform 1 0 308 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_449
timestamp 1554483974
transform 1 0 324 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_450
timestamp 1554483974
transform 1 0 332 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_399
timestamp 1554483974
transform 1 0 356 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_451
timestamp 1554483974
transform 1 0 388 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_414
timestamp 1554483974
transform 1 0 428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_415
timestamp 1554483974
transform 1 0 484 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_452
timestamp 1554483974
transform 1 0 404 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_362
timestamp 1554483974
transform 1 0 404 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_346
timestamp 1554483974
transform 1 0 524 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_453
timestamp 1554483974
transform 1 0 524 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_347
timestamp 1554483974
transform 1 0 564 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_416
timestamp 1554483974
transform 1 0 532 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_417
timestamp 1554483974
transform 1 0 548 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_418
timestamp 1554483974
transform 1 0 564 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_454
timestamp 1554483974
transform 1 0 540 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_455
timestamp 1554483974
transform 1 0 556 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_456
timestamp 1554483974
transform 1 0 604 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_341
timestamp 1554483974
transform 1 0 708 0 1 1035
box -3 -3 3 3
use M3_M2  M3_M2_348
timestamp 1554483974
transform 1 0 708 0 1 1025
box -3 -3 3 3
use M3_M2  M3_M2_342
timestamp 1554483974
transform 1 0 740 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_400
timestamp 1554483974
transform 1 0 724 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_349
timestamp 1554483974
transform 1 0 732 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_419
timestamp 1554483974
transform 1 0 644 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_420
timestamp 1554483974
transform 1 0 708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_421
timestamp 1554483974
transform 1 0 716 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_457
timestamp 1554483974
transform 1 0 620 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_458
timestamp 1554483974
transform 1 0 708 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_378
timestamp 1554483974
transform 1 0 620 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_422
timestamp 1554483974
transform 1 0 740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_459
timestamp 1554483974
transform 1 0 732 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_363
timestamp 1554483974
transform 1 0 732 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_364
timestamp 1554483974
transform 1 0 772 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_343
timestamp 1554483974
transform 1 0 836 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_423
timestamp 1554483974
transform 1 0 820 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_424
timestamp 1554483974
transform 1 0 868 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_425
timestamp 1554483974
transform 1 0 876 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_460
timestamp 1554483974
transform 1 0 788 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_461
timestamp 1554483974
transform 1 0 876 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_365
timestamp 1554483974
transform 1 0 876 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_379
timestamp 1554483974
transform 1 0 788 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_401
timestamp 1554483974
transform 1 0 900 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_462
timestamp 1554483974
transform 1 0 892 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_344
timestamp 1554483974
transform 1 0 916 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_402
timestamp 1554483974
transform 1 0 916 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_426
timestamp 1554483974
transform 1 0 924 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_463
timestamp 1554483974
transform 1 0 932 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_345
timestamp 1554483974
transform 1 0 980 0 1 1035
box -3 -3 3 3
use M2_M1  M2_M1_403
timestamp 1554483974
transform 1 0 980 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_464
timestamp 1554483974
transform 1 0 980 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_366
timestamp 1554483974
transform 1 0 964 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_367
timestamp 1554483974
transform 1 0 980 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_427
timestamp 1554483974
transform 1 0 1020 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_428
timestamp 1554483974
transform 1 0 1052 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_355
timestamp 1554483974
transform 1 0 1116 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_465
timestamp 1554483974
transform 1 0 1100 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_466
timestamp 1554483974
transform 1 0 1116 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_368
timestamp 1554483974
transform 1 0 1052 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_369
timestamp 1554483974
transform 1 0 1100 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_370
timestamp 1554483974
transform 1 0 1124 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_380
timestamp 1554483974
transform 1 0 1124 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_404
timestamp 1554483974
transform 1 0 1148 0 1 1025
box -2 -2 2 2
use M3_M2  M3_M2_350
timestamp 1554483974
transform 1 0 1156 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_405
timestamp 1554483974
transform 1 0 1180 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_429
timestamp 1554483974
transform 1 0 1156 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_430
timestamp 1554483974
transform 1 0 1172 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_356
timestamp 1554483974
transform 1 0 1180 0 1 1015
box -3 -3 3 3
use M3_M2  M3_M2_351
timestamp 1554483974
transform 1 0 1204 0 1 1025
box -3 -3 3 3
use M2_M1  M2_M1_431
timestamp 1554483974
transform 1 0 1196 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_467
timestamp 1554483974
transform 1 0 1172 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_468
timestamp 1554483974
transform 1 0 1180 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_432
timestamp 1554483974
transform 1 0 1220 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_433
timestamp 1554483974
transform 1 0 1252 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_469
timestamp 1554483974
transform 1 0 1212 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_371
timestamp 1554483974
transform 1 0 1212 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_470
timestamp 1554483974
transform 1 0 1300 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_381
timestamp 1554483974
transform 1 0 1300 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_434
timestamp 1554483974
transform 1 0 1316 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_471
timestamp 1554483974
transform 1 0 1324 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_372
timestamp 1554483974
transform 1 0 1324 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_472
timestamp 1554483974
transform 1 0 1356 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_373
timestamp 1554483974
transform 1 0 1348 0 1 995
box -3 -3 3 3
use M2_M1  M2_M1_406
timestamp 1554483974
transform 1 0 1364 0 1 1025
box -2 -2 2 2
use M2_M1  M2_M1_435
timestamp 1554483974
transform 1 0 1428 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_436
timestamp 1554483974
transform 1 0 1460 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_473
timestamp 1554483974
transform 1 0 1380 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_374
timestamp 1554483974
transform 1 0 1428 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_382
timestamp 1554483974
transform 1 0 1396 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_383
timestamp 1554483974
transform 1 0 1444 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_437
timestamp 1554483974
transform 1 0 1476 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_474
timestamp 1554483974
transform 1 0 1484 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_438
timestamp 1554483974
transform 1 0 1508 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_439
timestamp 1554483974
transform 1 0 1524 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_475
timestamp 1554483974
transform 1 0 1516 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_476
timestamp 1554483974
transform 1 0 1532 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_375
timestamp 1554483974
transform 1 0 1516 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_384
timestamp 1554483974
transform 1 0 1524 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_440
timestamp 1554483974
transform 1 0 1636 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_441
timestamp 1554483974
transform 1 0 1684 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_477
timestamp 1554483974
transform 1 0 1588 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_359
timestamp 1554483974
transform 1 0 1636 0 1 1005
box -3 -3 3 3
use M3_M2  M3_M2_360
timestamp 1554483974
transform 1 0 1668 0 1 1005
box -3 -3 3 3
use M2_M1  M2_M1_478
timestamp 1554483974
transform 1 0 1676 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_376
timestamp 1554483974
transform 1 0 1628 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_377
timestamp 1554483974
transform 1 0 1676 0 1 995
box -3 -3 3 3
use M3_M2  M3_M2_385
timestamp 1554483974
transform 1 0 1660 0 1 985
box -3 -3 3 3
use M3_M2  M3_M2_357
timestamp 1554483974
transform 1 0 1700 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_479
timestamp 1554483974
transform 1 0 1700 0 1 1005
box -2 -2 2 2
use M2_M1  M2_M1_442
timestamp 1554483974
transform 1 0 1708 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_443
timestamp 1554483974
transform 1 0 1724 0 1 1015
box -2 -2 2 2
use M3_M2  M3_M2_358
timestamp 1554483974
transform 1 0 1732 0 1 1015
box -3 -3 3 3
use M2_M1  M2_M1_444
timestamp 1554483974
transform 1 0 1740 0 1 1015
box -2 -2 2 2
use M2_M1  M2_M1_480
timestamp 1554483974
transform 1 0 1732 0 1 1005
box -2 -2 2 2
use M3_M2  M3_M2_386
timestamp 1554483974
transform 1 0 1740 0 1 985
box -3 -3 3 3
use M2_M1  M2_M1_481
timestamp 1554483974
transform 1 0 1756 0 1 1005
box -2 -2 2 2
use UART_VIA1  UART_VIA1_12
timestamp 1554483974
transform 1 0 48 0 1 970
box -10 -3 10 3
use FILL  FILL_411
timestamp 1554483974
transform 1 0 72 0 1 970
box -8 -3 16 105
use FILL  FILL_412
timestamp 1554483974
transform 1 0 80 0 1 970
box -8 -3 16 105
use FILL  FILL_413
timestamp 1554483974
transform 1 0 88 0 1 970
box -8 -3 16 105
use FILL  FILL_414
timestamp 1554483974
transform 1 0 96 0 1 970
box -8 -3 16 105
use NAND3X1  NAND3X1_4
timestamp 1554483974
transform -1 0 136 0 1 970
box -8 -3 40 105
use FILL  FILL_415
timestamp 1554483974
transform 1 0 136 0 1 970
box -8 -3 16 105
use FILL  FILL_416
timestamp 1554483974
transform 1 0 144 0 1 970
box -8 -3 16 105
use FILL  FILL_417
timestamp 1554483974
transform 1 0 152 0 1 970
box -8 -3 16 105
use OR2X1  OR2X1_1
timestamp 1554483974
transform 1 0 160 0 1 970
box -8 -3 40 105
use FILL  FILL_418
timestamp 1554483974
transform 1 0 192 0 1 970
box -8 -3 16 105
use FILL  FILL_419
timestamp 1554483974
transform 1 0 200 0 1 970
box -8 -3 16 105
use NOR2X1  NOR2X1_7
timestamp 1554483974
transform -1 0 232 0 1 970
box -8 -3 32 105
use INVX2  INVX2_22
timestamp 1554483974
transform 1 0 232 0 1 970
box -9 -3 26 105
use FILL  FILL_420
timestamp 1554483974
transform 1 0 248 0 1 970
box -8 -3 16 105
use FILL  FILL_421
timestamp 1554483974
transform 1 0 256 0 1 970
box -8 -3 16 105
use FILL  FILL_422
timestamp 1554483974
transform 1 0 264 0 1 970
box -8 -3 16 105
use FILL  FILL_431
timestamp 1554483974
transform 1 0 272 0 1 970
box -8 -3 16 105
use FILL  FILL_433
timestamp 1554483974
transform 1 0 280 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_8
timestamp 1554483974
transform -1 0 328 0 1 970
box -8 -3 46 105
use OAI21X1  OAI21X1_15
timestamp 1554483974
transform 1 0 328 0 1 970
box -8 -3 34 105
use FILL  FILL_434
timestamp 1554483974
transform 1 0 360 0 1 970
box -8 -3 16 105
use FILL  FILL_443
timestamp 1554483974
transform 1 0 368 0 1 970
box -8 -3 16 105
use FILL  FILL_445
timestamp 1554483974
transform 1 0 376 0 1 970
box -8 -3 16 105
use FILL  FILL_447
timestamp 1554483974
transform 1 0 384 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_18
timestamp 1554483974
transform 1 0 392 0 1 970
box -8 -3 104 105
use FILL  FILL_449
timestamp 1554483974
transform 1 0 488 0 1 970
box -8 -3 16 105
use FILL  FILL_456
timestamp 1554483974
transform 1 0 496 0 1 970
box -8 -3 16 105
use FILL  FILL_458
timestamp 1554483974
transform 1 0 504 0 1 970
box -8 -3 16 105
use FILL  FILL_460
timestamp 1554483974
transform 1 0 512 0 1 970
box -8 -3 16 105
use INVX2  INVX2_25
timestamp 1554483974
transform 1 0 520 0 1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_10
timestamp 1554483974
transform -1 0 576 0 1 970
box -8 -3 46 105
use FILL  FILL_462
timestamp 1554483974
transform 1 0 576 0 1 970
box -8 -3 16 105
use FILL  FILL_463
timestamp 1554483974
transform 1 0 584 0 1 970
box -8 -3 16 105
use FILL  FILL_464
timestamp 1554483974
transform 1 0 592 0 1 970
box -8 -3 16 105
use FILL  FILL_465
timestamp 1554483974
transform 1 0 600 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_19
timestamp 1554483974
transform 1 0 608 0 1 970
box -8 -3 104 105
use NAND2X1  NAND2X1_21
timestamp 1554483974
transform 1 0 704 0 1 970
box -8 -3 32 105
use INVX2  INVX2_26
timestamp 1554483974
transform 1 0 728 0 1 970
box -9 -3 26 105
use FILL  FILL_466
timestamp 1554483974
transform 1 0 744 0 1 970
box -8 -3 16 105
use FILL  FILL_467
timestamp 1554483974
transform 1 0 752 0 1 970
box -8 -3 16 105
use FILL  FILL_468
timestamp 1554483974
transform 1 0 760 0 1 970
box -8 -3 16 105
use FILL  FILL_469
timestamp 1554483974
transform 1 0 768 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_20
timestamp 1554483974
transform 1 0 776 0 1 970
box -8 -3 104 105
use NAND2X1  NAND2X1_22
timestamp 1554483974
transform 1 0 872 0 1 970
box -8 -3 32 105
use FILL  FILL_470
timestamp 1554483974
transform 1 0 896 0 1 970
box -8 -3 16 105
use FILL  FILL_487
timestamp 1554483974
transform 1 0 904 0 1 970
box -8 -3 16 105
use FILL  FILL_489
timestamp 1554483974
transform 1 0 912 0 1 970
box -8 -3 16 105
use FILL  FILL_491
timestamp 1554483974
transform 1 0 920 0 1 970
box -8 -3 16 105
use FILL  FILL_493
timestamp 1554483974
transform 1 0 928 0 1 970
box -8 -3 16 105
use FILL  FILL_495
timestamp 1554483974
transform 1 0 936 0 1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_19
timestamp 1554483974
transform 1 0 944 0 1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_25
timestamp 1554483974
transform -1 0 1000 0 1 970
box -8 -3 32 105
use FILL  FILL_497
timestamp 1554483974
transform 1 0 1000 0 1 970
box -8 -3 16 105
use FILL  FILL_498
timestamp 1554483974
transform 1 0 1008 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_22
timestamp 1554483974
transform -1 0 1112 0 1 970
box -8 -3 104 105
use INVX2  INVX2_28
timestamp 1554483974
transform 1 0 1112 0 1 970
box -9 -3 26 105
use FILL  FILL_499
timestamp 1554483974
transform 1 0 1128 0 1 970
box -8 -3 16 105
use FILL  FILL_500
timestamp 1554483974
transform 1 0 1136 0 1 970
box -8 -3 16 105
use FILL  FILL_501
timestamp 1554483974
transform 1 0 1144 0 1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_26
timestamp 1554483974
transform -1 0 1176 0 1 970
box -8 -3 32 105
use OAI21X1  OAI21X1_20
timestamp 1554483974
transform -1 0 1208 0 1 970
box -8 -3 34 105
use FILL  FILL_502
timestamp 1554483974
transform 1 0 1208 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_387
timestamp 1554483974
transform 1 0 1268 0 1 975
box -3 -3 3 3
use M3_M2  M3_M2_388
timestamp 1554483974
transform 1 0 1308 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_23
timestamp 1554483974
transform -1 0 1312 0 1 970
box -8 -3 104 105
use FILL  FILL_503
timestamp 1554483974
transform 1 0 1312 0 1 970
box -8 -3 16 105
use FILL  FILL_504
timestamp 1554483974
transform 1 0 1320 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_389
timestamp 1554483974
transform 1 0 1364 0 1 975
box -3 -3 3 3
use OAI21X1  OAI21X1_21
timestamp 1554483974
transform 1 0 1328 0 1 970
box -8 -3 34 105
use FILL  FILL_505
timestamp 1554483974
transform 1 0 1360 0 1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_24
timestamp 1554483974
transform 1 0 1368 0 1 970
box -8 -3 104 105
use FILL  FILL_506
timestamp 1554483974
transform 1 0 1464 0 1 970
box -8 -3 16 105
use FILL  FILL_507
timestamp 1554483974
transform 1 0 1472 0 1 970
box -8 -3 16 105
use FILL  FILL_508
timestamp 1554483974
transform 1 0 1480 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_390
timestamp 1554483974
transform 1 0 1500 0 1 975
box -3 -3 3 3
use FILL  FILL_509
timestamp 1554483974
transform 1 0 1488 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_391
timestamp 1554483974
transform 1 0 1532 0 1 975
box -3 -3 3 3
use OAI22X1  OAI22X1_11
timestamp 1554483974
transform -1 0 1536 0 1 970
box -8 -3 46 105
use FILL  FILL_510
timestamp 1554483974
transform 1 0 1536 0 1 970
box -8 -3 16 105
use FILL  FILL_511
timestamp 1554483974
transform 1 0 1544 0 1 970
box -8 -3 16 105
use FILL  FILL_512
timestamp 1554483974
transform 1 0 1552 0 1 970
box -8 -3 16 105
use FILL  FILL_513
timestamp 1554483974
transform 1 0 1560 0 1 970
box -8 -3 16 105
use FILL  FILL_514
timestamp 1554483974
transform 1 0 1568 0 1 970
box -8 -3 16 105
use M3_M2  M3_M2_392
timestamp 1554483974
transform 1 0 1588 0 1 975
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_25
timestamp 1554483974
transform 1 0 1576 0 1 970
box -8 -3 104 105
use M3_M2  M3_M2_393
timestamp 1554483974
transform 1 0 1692 0 1 975
box -3 -3 3 3
use INVX2  INVX2_29
timestamp 1554483974
transform 1 0 1672 0 1 970
box -9 -3 26 105
use FILL  FILL_515
timestamp 1554483974
transform 1 0 1688 0 1 970
box -8 -3 16 105
use FILL  FILL_530
timestamp 1554483974
transform 1 0 1696 0 1 970
box -8 -3 16 105
use FILL  FILL_532
timestamp 1554483974
transform 1 0 1704 0 1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_13
timestamp 1554483974
transform -1 0 1752 0 1 970
box -8 -3 46 105
use FILL  FILL_533
timestamp 1554483974
transform 1 0 1752 0 1 970
box -8 -3 16 105
use FILL  FILL_534
timestamp 1554483974
transform 1 0 1760 0 1 970
box -8 -3 16 105
use FILL  FILL_541
timestamp 1554483974
transform 1 0 1768 0 1 970
box -8 -3 16 105
use UART_VIA1  UART_VIA1_13
timestamp 1554483974
transform 1 0 1801 0 1 970
box -10 -3 10 3
use M3_M2  M3_M2_414
timestamp 1554483974
transform 1 0 68 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_485
timestamp 1554483974
transform 1 0 156 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_522
timestamp 1554483974
transform 1 0 68 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_523
timestamp 1554483974
transform 1 0 132 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_486
timestamp 1554483974
transform 1 0 180 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_524
timestamp 1554483974
transform 1 0 172 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_415
timestamp 1554483974
transform 1 0 188 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_558
timestamp 1554483974
transform 1 0 196 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_525
timestamp 1554483974
transform 1 0 212 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_422
timestamp 1554483974
transform 1 0 228 0 1 925
box -3 -3 3 3
use M3_M2  M3_M2_399
timestamp 1554483974
transform 1 0 252 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_487
timestamp 1554483974
transform 1 0 252 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_400
timestamp 1554483974
transform 1 0 316 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_488
timestamp 1554483974
transform 1 0 340 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_423
timestamp 1554483974
transform 1 0 340 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_526
timestamp 1554483974
transform 1 0 356 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_428
timestamp 1554483974
transform 1 0 356 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_416
timestamp 1554483974
transform 1 0 388 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_559
timestamp 1554483974
transform 1 0 380 0 1 915
box -2 -2 2 2
use M2_M1  M2_M1_489
timestamp 1554483974
transform 1 0 404 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_417
timestamp 1554483974
transform 1 0 412 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_490
timestamp 1554483974
transform 1 0 420 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_527
timestamp 1554483974
transform 1 0 412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_528
timestamp 1554483974
transform 1 0 428 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_529
timestamp 1554483974
transform 1 0 452 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_429
timestamp 1554483974
transform 1 0 428 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_491
timestamp 1554483974
transform 1 0 484 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_394
timestamp 1554483974
transform 1 0 604 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_395
timestamp 1554483974
transform 1 0 628 0 1 965
box -3 -3 3 3
use M3_M2  M3_M2_401
timestamp 1554483974
transform 1 0 532 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_402
timestamp 1554483974
transform 1 0 620 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_492
timestamp 1554483974
transform 1 0 532 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_530
timestamp 1554483974
transform 1 0 556 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_531
timestamp 1554483974
transform 1 0 628 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_430
timestamp 1554483974
transform 1 0 628 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_493
timestamp 1554483974
transform 1 0 684 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_403
timestamp 1554483974
transform 1 0 740 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_494
timestamp 1554483974
transform 1 0 732 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_495
timestamp 1554483974
transform 1 0 740 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_532
timestamp 1554483974
transform 1 0 716 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_533
timestamp 1554483974
transform 1 0 724 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_560
timestamp 1554483974
transform 1 0 700 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_431
timestamp 1554483974
transform 1 0 724 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_496
timestamp 1554483974
transform 1 0 764 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_561
timestamp 1554483974
transform 1 0 772 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_437
timestamp 1554483974
transform 1 0 772 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_404
timestamp 1554483974
transform 1 0 796 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_497
timestamp 1554483974
transform 1 0 796 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_534
timestamp 1554483974
transform 1 0 812 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_535
timestamp 1554483974
transform 1 0 836 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_498
timestamp 1554483974
transform 1 0 868 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_405
timestamp 1554483974
transform 1 0 892 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_562
timestamp 1554483974
transform 1 0 876 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_438
timestamp 1554483974
transform 1 0 876 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_499
timestamp 1554483974
transform 1 0 908 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_439
timestamp 1554483974
transform 1 0 900 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_500
timestamp 1554483974
transform 1 0 932 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_406
timestamp 1554483974
transform 1 0 956 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_501
timestamp 1554483974
transform 1 0 956 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_536
timestamp 1554483974
transform 1 0 964 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_432
timestamp 1554483974
transform 1 0 964 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_407
timestamp 1554483974
transform 1 0 988 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_502
timestamp 1554483974
transform 1 0 988 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_537
timestamp 1554483974
transform 1 0 996 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_424
timestamp 1554483974
transform 1 0 1004 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_503
timestamp 1554483974
transform 1 0 1036 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_538
timestamp 1554483974
transform 1 0 1012 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_539
timestamp 1554483974
transform 1 0 1028 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_540
timestamp 1554483974
transform 1 0 1044 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_433
timestamp 1554483974
transform 1 0 1012 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_434
timestamp 1554483974
transform 1 0 1044 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_440
timestamp 1554483974
transform 1 0 1028 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_444
timestamp 1554483974
transform 1 0 1044 0 1 895
box -3 -3 3 3
use M2_M1  M2_M1_504
timestamp 1554483974
transform 1 0 1068 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_445
timestamp 1554483974
transform 1 0 1068 0 1 895
box -3 -3 3 3
use M3_M2  M3_M2_418
timestamp 1554483974
transform 1 0 1100 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_541
timestamp 1554483974
transform 1 0 1092 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_542
timestamp 1554483974
transform 1 0 1100 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_396
timestamp 1554483974
transform 1 0 1172 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_397
timestamp 1554483974
transform 1 0 1204 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_398
timestamp 1554483974
transform 1 0 1260 0 1 955
box -3 -3 3 3
use M3_M2  M3_M2_408
timestamp 1554483974
transform 1 0 1236 0 1 945
box -3 -3 3 3
use M3_M2  M3_M2_409
timestamp 1554483974
transform 1 0 1252 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_505
timestamp 1554483974
transform 1 0 1124 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_506
timestamp 1554483974
transform 1 0 1212 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_419
timestamp 1554483974
transform 1 0 1220 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_543
timestamp 1554483974
transform 1 0 1172 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_544
timestamp 1554483974
transform 1 0 1204 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_545
timestamp 1554483974
transform 1 0 1212 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_546
timestamp 1554483974
transform 1 0 1220 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_547
timestamp 1554483974
transform 1 0 1236 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_563
timestamp 1554483974
transform 1 0 1108 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_435
timestamp 1554483974
transform 1 0 1196 0 1 915
box -3 -3 3 3
use M3_M2  M3_M2_436
timestamp 1554483974
transform 1 0 1220 0 1 915
box -3 -3 3 3
use M2_M1  M2_M1_507
timestamp 1554483974
transform 1 0 1244 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_508
timestamp 1554483974
transform 1 0 1260 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_564
timestamp 1554483974
transform 1 0 1244 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_410
timestamp 1554483974
transform 1 0 1348 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_509
timestamp 1554483974
transform 1 0 1308 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_411
timestamp 1554483974
transform 1 0 1412 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_510
timestamp 1554483974
transform 1 0 1364 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_511
timestamp 1554483974
transform 1 0 1412 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_548
timestamp 1554483974
transform 1 0 1348 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_565
timestamp 1554483974
transform 1 0 1316 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_441
timestamp 1554483974
transform 1 0 1316 0 1 905
box -3 -3 3 3
use M3_M2  M3_M2_425
timestamp 1554483974
transform 1 0 1372 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_549
timestamp 1554483974
transform 1 0 1412 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_566
timestamp 1554483974
transform 1 0 1372 0 1 915
box -2 -2 2 2
use M3_M2  M3_M2_442
timestamp 1554483974
transform 1 0 1412 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_512
timestamp 1554483974
transform 1 0 1460 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_513
timestamp 1554483974
transform 1 0 1476 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_412
timestamp 1554483974
transform 1 0 1492 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_550
timestamp 1554483974
transform 1 0 1484 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_413
timestamp 1554483974
transform 1 0 1508 0 1 945
box -3 -3 3 3
use M2_M1  M2_M1_514
timestamp 1554483974
transform 1 0 1508 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_515
timestamp 1554483974
transform 1 0 1516 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_551
timestamp 1554483974
transform 1 0 1500 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_552
timestamp 1554483974
transform 1 0 1508 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_443
timestamp 1554483974
transform 1 0 1516 0 1 905
box -3 -3 3 3
use M2_M1  M2_M1_516
timestamp 1554483974
transform 1 0 1564 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_553
timestamp 1554483974
transform 1 0 1572 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_554
timestamp 1554483974
transform 1 0 1596 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_517
timestamp 1554483974
transform 1 0 1628 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_518
timestamp 1554483974
transform 1 0 1636 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_420
timestamp 1554483974
transform 1 0 1644 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_519
timestamp 1554483974
transform 1 0 1668 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_421
timestamp 1554483974
transform 1 0 1676 0 1 935
box -3 -3 3 3
use M2_M1  M2_M1_520
timestamp 1554483974
transform 1 0 1684 0 1 935
box -2 -2 2 2
use M3_M2  M3_M2_426
timestamp 1554483974
transform 1 0 1652 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_555
timestamp 1554483974
transform 1 0 1660 0 1 925
box -2 -2 2 2
use M2_M1  M2_M1_556
timestamp 1554483974
transform 1 0 1676 0 1 925
box -2 -2 2 2
use M3_M2  M3_M2_427
timestamp 1554483974
transform 1 0 1700 0 1 925
box -3 -3 3 3
use M2_M1  M2_M1_521
timestamp 1554483974
transform 1 0 1724 0 1 935
box -2 -2 2 2
use M2_M1  M2_M1_557
timestamp 1554483974
transform 1 0 1756 0 1 925
box -2 -2 2 2
use UART_VIA1  UART_VIA1_14
timestamp 1554483974
transform 1 0 24 0 1 870
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_17
timestamp 1554483974
transform -1 0 168 0 -1 970
box -8 -3 104 105
use FILL  FILL_423
timestamp 1554483974
transform 1 0 168 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_19
timestamp 1554483974
transform 1 0 176 0 -1 970
box -8 -3 32 105
use FILL  FILL_424
timestamp 1554483974
transform 1 0 200 0 -1 970
box -8 -3 16 105
use FILL  FILL_425
timestamp 1554483974
transform 1 0 208 0 -1 970
box -8 -3 16 105
use FILL  FILL_426
timestamp 1554483974
transform 1 0 216 0 -1 970
box -8 -3 16 105
use FILL  FILL_427
timestamp 1554483974
transform 1 0 224 0 -1 970
box -8 -3 16 105
use FILL  FILL_428
timestamp 1554483974
transform 1 0 232 0 -1 970
box -8 -3 16 105
use FILL  FILL_429
timestamp 1554483974
transform 1 0 240 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_23
timestamp 1554483974
transform 1 0 248 0 -1 970
box -9 -3 26 105
use FILL  FILL_430
timestamp 1554483974
transform 1 0 264 0 -1 970
box -8 -3 16 105
use FILL  FILL_432
timestamp 1554483974
transform 1 0 272 0 -1 970
box -8 -3 16 105
use FILL  FILL_435
timestamp 1554483974
transform 1 0 280 0 -1 970
box -8 -3 16 105
use FILL  FILL_436
timestamp 1554483974
transform 1 0 288 0 -1 970
box -8 -3 16 105
use FILL  FILL_437
timestamp 1554483974
transform 1 0 296 0 -1 970
box -8 -3 16 105
use FILL  FILL_438
timestamp 1554483974
transform 1 0 304 0 -1 970
box -8 -3 16 105
use FILL  FILL_439
timestamp 1554483974
transform 1 0 312 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_20
timestamp 1554483974
transform 1 0 320 0 -1 970
box -8 -3 32 105
use FILL  FILL_440
timestamp 1554483974
transform 1 0 344 0 -1 970
box -8 -3 16 105
use FILL  FILL_441
timestamp 1554483974
transform 1 0 352 0 -1 970
box -8 -3 16 105
use FILL  FILL_442
timestamp 1554483974
transform 1 0 360 0 -1 970
box -8 -3 16 105
use FILL  FILL_444
timestamp 1554483974
transform 1 0 368 0 -1 970
box -8 -3 16 105
use FILL  FILL_446
timestamp 1554483974
transform 1 0 376 0 -1 970
box -8 -3 16 105
use FILL  FILL_448
timestamp 1554483974
transform 1 0 384 0 -1 970
box -8 -3 16 105
use FILL  FILL_450
timestamp 1554483974
transform 1 0 392 0 -1 970
box -8 -3 16 105
use OAI22X1  OAI22X1_9
timestamp 1554483974
transform -1 0 440 0 -1 970
box -8 -3 46 105
use INVX2  INVX2_24
timestamp 1554483974
transform -1 0 456 0 -1 970
box -9 -3 26 105
use FILL  FILL_451
timestamp 1554483974
transform 1 0 456 0 -1 970
box -8 -3 16 105
use FILL  FILL_452
timestamp 1554483974
transform 1 0 464 0 -1 970
box -8 -3 16 105
use FILL  FILL_453
timestamp 1554483974
transform 1 0 472 0 -1 970
box -8 -3 16 105
use FILL  FILL_454
timestamp 1554483974
transform 1 0 480 0 -1 970
box -8 -3 16 105
use FILL  FILL_455
timestamp 1554483974
transform 1 0 488 0 -1 970
box -8 -3 16 105
use FILL  FILL_457
timestamp 1554483974
transform 1 0 496 0 -1 970
box -8 -3 16 105
use FILL  FILL_459
timestamp 1554483974
transform 1 0 504 0 -1 970
box -8 -3 16 105
use FILL  FILL_461
timestamp 1554483974
transform 1 0 512 0 -1 970
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_21
timestamp 1554483974
transform 1 0 520 0 -1 970
box -8 -3 104 105
use INVX2  INVX2_27
timestamp 1554483974
transform 1 0 616 0 -1 970
box -9 -3 26 105
use FILL  FILL_471
timestamp 1554483974
transform 1 0 632 0 -1 970
box -8 -3 16 105
use FILL  FILL_472
timestamp 1554483974
transform 1 0 640 0 -1 970
box -8 -3 16 105
use FILL  FILL_473
timestamp 1554483974
transform 1 0 648 0 -1 970
box -8 -3 16 105
use FILL  FILL_474
timestamp 1554483974
transform 1 0 656 0 -1 970
box -8 -3 16 105
use FILL  FILL_475
timestamp 1554483974
transform 1 0 664 0 -1 970
box -8 -3 16 105
use FILL  FILL_476
timestamp 1554483974
transform 1 0 672 0 -1 970
box -8 -3 16 105
use FILL  FILL_477
timestamp 1554483974
transform 1 0 680 0 -1 970
box -8 -3 16 105
use FILL  FILL_478
timestamp 1554483974
transform 1 0 688 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_16
timestamp 1554483974
transform -1 0 728 0 -1 970
box -8 -3 34 105
use FILL  FILL_479
timestamp 1554483974
transform 1 0 728 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_17
timestamp 1554483974
transform 1 0 736 0 -1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_23
timestamp 1554483974
transform -1 0 792 0 -1 970
box -8 -3 32 105
use FILL  FILL_480
timestamp 1554483974
transform 1 0 792 0 -1 970
box -8 -3 16 105
use FILL  FILL_481
timestamp 1554483974
transform 1 0 800 0 -1 970
box -8 -3 16 105
use FILL  FILL_482
timestamp 1554483974
transform 1 0 808 0 -1 970
box -8 -3 16 105
use FILL  FILL_483
timestamp 1554483974
transform 1 0 816 0 -1 970
box -8 -3 16 105
use FILL  FILL_484
timestamp 1554483974
transform 1 0 824 0 -1 970
box -8 -3 16 105
use FILL  FILL_485
timestamp 1554483974
transform 1 0 832 0 -1 970
box -8 -3 16 105
use OAI21X1  OAI21X1_18
timestamp 1554483974
transform 1 0 840 0 -1 970
box -8 -3 34 105
use NAND2X1  NAND2X1_24
timestamp 1554483974
transform -1 0 896 0 -1 970
box -8 -3 32 105
use FILL  FILL_486
timestamp 1554483974
transform 1 0 896 0 -1 970
box -8 -3 16 105
use FILL  FILL_488
timestamp 1554483974
transform 1 0 904 0 -1 970
box -8 -3 16 105
use FILL  FILL_490
timestamp 1554483974
transform 1 0 912 0 -1 970
box -8 -3 16 105
use FILL  FILL_492
timestamp 1554483974
transform 1 0 920 0 -1 970
box -8 -3 16 105
use FILL  FILL_494
timestamp 1554483974
transform 1 0 928 0 -1 970
box -8 -3 16 105
use FILL  FILL_496
timestamp 1554483974
transform 1 0 936 0 -1 970
box -8 -3 16 105
use FILL  FILL_516
timestamp 1554483974
transform 1 0 944 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_8
timestamp 1554483974
transform 1 0 952 0 -1 970
box -8 -3 40 105
use FILL  FILL_517
timestamp 1554483974
transform 1 0 984 0 -1 970
box -8 -3 16 105
use FILL  FILL_518
timestamp 1554483974
transform 1 0 992 0 -1 970
box -8 -3 16 105
use AND2X2  AND2X2_9
timestamp 1554483974
transform 1 0 1000 0 -1 970
box -8 -3 40 105
use AND2X2  AND2X2_10
timestamp 1554483974
transform 1 0 1032 0 -1 970
box -8 -3 40 105
use FILL  FILL_519
timestamp 1554483974
transform 1 0 1064 0 -1 970
box -8 -3 16 105
use FILL  FILL_520
timestamp 1554483974
transform 1 0 1072 0 -1 970
box -8 -3 16 105
use FILL  FILL_521
timestamp 1554483974
transform 1 0 1080 0 -1 970
box -8 -3 16 105
use NAND2X1  NAND2X1_27
timestamp 1554483974
transform 1 0 1088 0 -1 970
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_26
timestamp 1554483974
transform 1 0 1112 0 -1 970
box -8 -3 104 105
use OAI21X1  OAI21X1_22
timestamp 1554483974
transform 1 0 1208 0 -1 970
box -8 -3 34 105
use FILL  FILL_522
timestamp 1554483974
transform 1 0 1240 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_30
timestamp 1554483974
transform -1 0 1264 0 -1 970
box -9 -3 26 105
use FILL  FILL_523
timestamp 1554483974
transform 1 0 1264 0 -1 970
box -8 -3 16 105
use FILL  FILL_524
timestamp 1554483974
transform 1 0 1272 0 -1 970
box -8 -3 16 105
use FILL  FILL_525
timestamp 1554483974
transform 1 0 1280 0 -1 970
box -8 -3 16 105
use FILL  FILL_526
timestamp 1554483974
transform 1 0 1288 0 -1 970
box -8 -3 16 105
use LATCH  LATCH_8
timestamp 1554483974
transform 1 0 1296 0 -1 970
box -8 -3 64 105
use LATCH  LATCH_9
timestamp 1554483974
transform 1 0 1352 0 -1 970
box -8 -3 64 105
use XOR2X1  XOR2X1_9
timestamp 1554483974
transform 1 0 1408 0 -1 970
box -8 -3 64 105
use NOR2X1  NOR2X1_8
timestamp 1554483974
transform 1 0 1464 0 -1 970
box -8 -3 32 105
use FILL  FILL_527
timestamp 1554483974
transform 1 0 1488 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_31
timestamp 1554483974
transform -1 0 1512 0 -1 970
box -9 -3 26 105
use M3_M2  M3_M2_446
timestamp 1554483974
transform 1 0 1548 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_10
timestamp 1554483974
transform -1 0 1568 0 -1 970
box -8 -3 64 105
use M3_M2  M3_M2_447
timestamp 1554483974
transform 1 0 1596 0 1 875
box -3 -3 3 3
use XOR2X1  XOR2X1_11
timestamp 1554483974
transform 1 0 1568 0 -1 970
box -8 -3 64 105
use FILL  FILL_528
timestamp 1554483974
transform 1 0 1624 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_32
timestamp 1554483974
transform 1 0 1632 0 -1 970
box -9 -3 26 105
use OAI22X1  OAI22X1_12
timestamp 1554483974
transform 1 0 1648 0 -1 970
box -8 -3 46 105
use FILL  FILL_529
timestamp 1554483974
transform 1 0 1688 0 -1 970
box -8 -3 16 105
use FILL  FILL_531
timestamp 1554483974
transform 1 0 1696 0 -1 970
box -8 -3 16 105
use FILL  FILL_535
timestamp 1554483974
transform 1 0 1704 0 -1 970
box -8 -3 16 105
use FILL  FILL_536
timestamp 1554483974
transform 1 0 1712 0 -1 970
box -8 -3 16 105
use FILL  FILL_537
timestamp 1554483974
transform 1 0 1720 0 -1 970
box -8 -3 16 105
use FILL  FILL_538
timestamp 1554483974
transform 1 0 1728 0 -1 970
box -8 -3 16 105
use FILL  FILL_539
timestamp 1554483974
transform 1 0 1736 0 -1 970
box -8 -3 16 105
use INVX2  INVX2_33
timestamp 1554483974
transform 1 0 1744 0 -1 970
box -9 -3 26 105
use FILL  FILL_540
timestamp 1554483974
transform 1 0 1760 0 -1 970
box -8 -3 16 105
use FILL  FILL_542
timestamp 1554483974
transform 1 0 1768 0 -1 970
box -8 -3 16 105
use UART_VIA1  UART_VIA1_15
timestamp 1554483974
transform 1 0 1825 0 1 870
box -10 -3 10 3
use M3_M2  M3_M2_448
timestamp 1554483974
transform 1 0 68 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_468
timestamp 1554483974
transform 1 0 68 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_469
timestamp 1554483974
transform 1 0 84 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_572
timestamp 1554483974
transform 1 0 108 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_470
timestamp 1554483974
transform 1 0 124 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_588
timestamp 1554483974
transform 1 0 124 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_589
timestamp 1554483974
transform 1 0 132 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_621
timestamp 1554483974
transform 1 0 108 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_622
timestamp 1554483974
transform 1 0 140 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_488
timestamp 1554483974
transform 1 0 140 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_462
timestamp 1554483974
transform 1 0 188 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_573
timestamp 1554483974
transform 1 0 172 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_590
timestamp 1554483974
transform 1 0 188 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_591
timestamp 1554483974
transform 1 0 196 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_592
timestamp 1554483974
transform 1 0 204 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_489
timestamp 1554483974
transform 1 0 204 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_623
timestamp 1554483974
transform 1 0 228 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_463
timestamp 1554483974
transform 1 0 260 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_574
timestamp 1554483974
transform 1 0 260 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_593
timestamp 1554483974
transform 1 0 252 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_575
timestamp 1554483974
transform 1 0 292 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_452
timestamp 1554483974
transform 1 0 340 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_567
timestamp 1554483974
transform 1 0 324 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_471
timestamp 1554483974
transform 1 0 324 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_568
timestamp 1554483974
transform 1 0 348 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_569
timestamp 1554483974
transform 1 0 356 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_576
timestamp 1554483974
transform 1 0 340 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_594
timestamp 1554483974
transform 1 0 324 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_595
timestamp 1554483974
transform 1 0 348 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_453
timestamp 1554483974
transform 1 0 436 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_570
timestamp 1554483974
transform 1 0 420 0 1 835
box -2 -2 2 2
use M2_M1  M2_M1_577
timestamp 1554483974
transform 1 0 404 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_578
timestamp 1554483974
transform 1 0 412 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_472
timestamp 1554483974
transform 1 0 428 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_579
timestamp 1554483974
transform 1 0 436 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_596
timestamp 1554483974
transform 1 0 428 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_597
timestamp 1554483974
transform 1 0 452 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_624
timestamp 1554483974
transform 1 0 476 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_449
timestamp 1554483974
transform 1 0 532 0 1 865
box -3 -3 3 3
use M3_M2  M3_M2_473
timestamp 1554483974
transform 1 0 540 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_625
timestamp 1554483974
transform 1 0 540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_626
timestamp 1554483974
transform 1 0 548 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_498
timestamp 1554483974
transform 1 0 548 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_454
timestamp 1554483974
transform 1 0 564 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_580
timestamp 1554483974
transform 1 0 564 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_474
timestamp 1554483974
transform 1 0 620 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_598
timestamp 1554483974
transform 1 0 620 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_599
timestamp 1554483974
transform 1 0 676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_627
timestamp 1554483974
transform 1 0 596 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_499
timestamp 1554483974
transform 1 0 676 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_455
timestamp 1554483974
transform 1 0 772 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_600
timestamp 1554483974
transform 1 0 756 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_601
timestamp 1554483974
transform 1 0 812 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_628
timestamp 1554483974
transform 1 0 732 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_490
timestamp 1554483974
transform 1 0 812 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_602
timestamp 1554483974
transform 1 0 868 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_629
timestamp 1554483974
transform 1 0 844 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_603
timestamp 1554483974
transform 1 0 932 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_486
timestamp 1554483974
transform 1 0 932 0 1 805
box -3 -3 3 3
use M2_M1  M2_M1_630
timestamp 1554483974
transform 1 0 948 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_475
timestamp 1554483974
transform 1 0 964 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_604
timestamp 1554483974
transform 1 0 964 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_500
timestamp 1554483974
transform 1 0 956 0 1 785
box -3 -3 3 3
use M2_M1  M2_M1_631
timestamp 1554483974
transform 1 0 988 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_487
timestamp 1554483974
transform 1 0 996 0 1 805
box -3 -3 3 3
use M3_M2  M3_M2_491
timestamp 1554483974
transform 1 0 988 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_464
timestamp 1554483974
transform 1 0 1012 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_605
timestamp 1554483974
transform 1 0 1012 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_476
timestamp 1554483974
transform 1 0 1028 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_606
timestamp 1554483974
transform 1 0 1028 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_456
timestamp 1554483974
transform 1 0 1068 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_607
timestamp 1554483974
transform 1 0 1068 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_450
timestamp 1554483974
transform 1 0 1092 0 1 855
box -3 -3 3 3
use M3_M2  M3_M2_465
timestamp 1554483974
transform 1 0 1092 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_581
timestamp 1554483974
transform 1 0 1092 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_632
timestamp 1554483974
transform 1 0 1084 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_492
timestamp 1554483974
transform 1 0 1084 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_582
timestamp 1554483974
transform 1 0 1148 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_477
timestamp 1554483974
transform 1 0 1164 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_633
timestamp 1554483974
transform 1 0 1172 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_608
timestamp 1554483974
transform 1 0 1180 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_609
timestamp 1554483974
transform 1 0 1212 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_634
timestamp 1554483974
transform 1 0 1212 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_457
timestamp 1554483974
transform 1 0 1276 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_583
timestamp 1554483974
transform 1 0 1276 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_635
timestamp 1554483974
transform 1 0 1268 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_493
timestamp 1554483974
transform 1 0 1268 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_610
timestamp 1554483974
transform 1 0 1332 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_494
timestamp 1554483974
transform 1 0 1324 0 1 795
box -3 -3 3 3
use M3_M2  M3_M2_501
timestamp 1554483974
transform 1 0 1332 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_451
timestamp 1554483974
transform 1 0 1356 0 1 855
box -3 -3 3 3
use M2_M1  M2_M1_584
timestamp 1554483974
transform 1 0 1356 0 1 825
box -2 -2 2 2
use M3_M2  M3_M2_481
timestamp 1554483974
transform 1 0 1348 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_482
timestamp 1554483974
transform 1 0 1372 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_636
timestamp 1554483974
transform 1 0 1348 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_495
timestamp 1554483974
transform 1 0 1348 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_637
timestamp 1554483974
transform 1 0 1412 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_585
timestamp 1554483974
transform 1 0 1476 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_638
timestamp 1554483974
transform 1 0 1468 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_611
timestamp 1554483974
transform 1 0 1484 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_458
timestamp 1554483974
transform 1 0 1508 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_571
timestamp 1554483974
transform 1 0 1508 0 1 835
box -2 -2 2 2
use M3_M2  M3_M2_478
timestamp 1554483974
transform 1 0 1508 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_459
timestamp 1554483974
transform 1 0 1532 0 1 845
box -3 -3 3 3
use M2_M1  M2_M1_586
timestamp 1554483974
transform 1 0 1516 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_612
timestamp 1554483974
transform 1 0 1500 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_613
timestamp 1554483974
transform 1 0 1548 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_483
timestamp 1554483974
transform 1 0 1572 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_466
timestamp 1554483974
transform 1 0 1604 0 1 835
box -3 -3 3 3
use M2_M1  M2_M1_614
timestamp 1554483974
transform 1 0 1596 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_639
timestamp 1554483974
transform 1 0 1532 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_640
timestamp 1554483974
transform 1 0 1540 0 1 805
box -2 -2 2 2
use M2_M1  M2_M1_643
timestamp 1554483974
transform 1 0 1524 0 1 795
box -2 -2 2 2
use M3_M2  M3_M2_502
timestamp 1554483974
transform 1 0 1564 0 1 785
box -3 -3 3 3
use M3_M2  M3_M2_460
timestamp 1554483974
transform 1 0 1644 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_461
timestamp 1554483974
transform 1 0 1676 0 1 845
box -3 -3 3 3
use M3_M2  M3_M2_467
timestamp 1554483974
transform 1 0 1660 0 1 835
box -3 -3 3 3
use M3_M2  M3_M2_479
timestamp 1554483974
transform 1 0 1636 0 1 825
box -3 -3 3 3
use M3_M2  M3_M2_484
timestamp 1554483974
transform 1 0 1628 0 1 815
box -3 -3 3 3
use M2_M1  M2_M1_587
timestamp 1554483974
transform 1 0 1676 0 1 825
box -2 -2 2 2
use M2_M1  M2_M1_615
timestamp 1554483974
transform 1 0 1636 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_616
timestamp 1554483974
transform 1 0 1652 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_617
timestamp 1554483974
transform 1 0 1660 0 1 815
box -2 -2 2 2
use M3_M2  M3_M2_485
timestamp 1554483974
transform 1 0 1668 0 1 815
box -3 -3 3 3
use M3_M2  M3_M2_480
timestamp 1554483974
transform 1 0 1772 0 1 825
box -3 -3 3 3
use M2_M1  M2_M1_618
timestamp 1554483974
transform 1 0 1676 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_619
timestamp 1554483974
transform 1 0 1732 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_620
timestamp 1554483974
transform 1 0 1772 0 1 815
box -2 -2 2 2
use M2_M1  M2_M1_641
timestamp 1554483974
transform 1 0 1652 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_496
timestamp 1554483974
transform 1 0 1652 0 1 795
box -3 -3 3 3
use M2_M1  M2_M1_642
timestamp 1554483974
transform 1 0 1692 0 1 805
box -2 -2 2 2
use M3_M2  M3_M2_497
timestamp 1554483974
transform 1 0 1724 0 1 795
box -3 -3 3 3
use UART_VIA1  UART_VIA1_16
timestamp 1554483974
transform 1 0 48 0 1 770
box -10 -3 10 3
use FILL  FILL_543
timestamp 1554483974
transform 1 0 72 0 1 770
box -8 -3 16 105
use FILL  FILL_544
timestamp 1554483974
transform 1 0 80 0 1 770
box -8 -3 16 105
use FILL  FILL_545
timestamp 1554483974
transform 1 0 88 0 1 770
box -8 -3 16 105
use FILL  FILL_546
timestamp 1554483974
transform 1 0 96 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_23
timestamp 1554483974
transform -1 0 136 0 1 770
box -8 -3 34 105
use FILL  FILL_547
timestamp 1554483974
transform 1 0 136 0 1 770
box -8 -3 16 105
use FILL  FILL_548
timestamp 1554483974
transform 1 0 144 0 1 770
box -8 -3 16 105
use FILL  FILL_549
timestamp 1554483974
transform 1 0 152 0 1 770
box -8 -3 16 105
use FILL  FILL_550
timestamp 1554483974
transform 1 0 160 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_24
timestamp 1554483974
transform -1 0 200 0 1 770
box -8 -3 34 105
use FILL  FILL_551
timestamp 1554483974
transform 1 0 200 0 1 770
box -8 -3 16 105
use FILL  FILL_552
timestamp 1554483974
transform 1 0 208 0 1 770
box -8 -3 16 105
use FILL  FILL_553
timestamp 1554483974
transform 1 0 216 0 1 770
box -8 -3 16 105
use FILL  FILL_554
timestamp 1554483974
transform 1 0 224 0 1 770
box -8 -3 16 105
use FILL  FILL_555
timestamp 1554483974
transform 1 0 232 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_28
timestamp 1554483974
transform 1 0 240 0 1 770
box -8 -3 32 105
use FILL  FILL_556
timestamp 1554483974
transform 1 0 264 0 1 770
box -8 -3 16 105
use FILL  FILL_557
timestamp 1554483974
transform 1 0 272 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_503
timestamp 1554483974
transform 1 0 292 0 1 775
box -3 -3 3 3
use FILL  FILL_558
timestamp 1554483974
transform 1 0 280 0 1 770
box -8 -3 16 105
use FILL  FILL_559
timestamp 1554483974
transform 1 0 288 0 1 770
box -8 -3 16 105
use FILL  FILL_560
timestamp 1554483974
transform 1 0 296 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_5
timestamp 1554483974
transform -1 0 336 0 1 770
box -8 -3 40 105
use NAND3X1  NAND3X1_6
timestamp 1554483974
transform 1 0 336 0 1 770
box -8 -3 40 105
use FILL  FILL_561
timestamp 1554483974
transform 1 0 368 0 1 770
box -8 -3 16 105
use FILL  FILL_568
timestamp 1554483974
transform 1 0 376 0 1 770
box -8 -3 16 105
use FILL  FILL_570
timestamp 1554483974
transform 1 0 384 0 1 770
box -8 -3 16 105
use FILL  FILL_572
timestamp 1554483974
transform 1 0 392 0 1 770
box -8 -3 16 105
use FILL  FILL_574
timestamp 1554483974
transform 1 0 400 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_504
timestamp 1554483974
transform 1 0 444 0 1 775
box -3 -3 3 3
use NAND3X1  NAND3X1_8
timestamp 1554483974
transform -1 0 440 0 1 770
box -8 -3 40 105
use FILL  FILL_575
timestamp 1554483974
transform 1 0 440 0 1 770
box -8 -3 16 105
use FILL  FILL_576
timestamp 1554483974
transform 1 0 448 0 1 770
box -8 -3 16 105
use FILL  FILL_581
timestamp 1554483974
transform 1 0 456 0 1 770
box -8 -3 16 105
use FILL  FILL_583
timestamp 1554483974
transform 1 0 464 0 1 770
box -8 -3 16 105
use FILL  FILL_585
timestamp 1554483974
transform 1 0 472 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_25
timestamp 1554483974
transform 1 0 480 0 1 770
box -8 -3 34 105
use FILL  FILL_587
timestamp 1554483974
transform 1 0 512 0 1 770
box -8 -3 16 105
use FILL  FILL_591
timestamp 1554483974
transform 1 0 520 0 1 770
box -8 -3 16 105
use FILL  FILL_593
timestamp 1554483974
transform 1 0 528 0 1 770
box -8 -3 16 105
use FILL  FILL_594
timestamp 1554483974
transform 1 0 536 0 1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_30
timestamp 1554483974
transform 1 0 544 0 1 770
box -8 -3 32 105
use FILL  FILL_595
timestamp 1554483974
transform 1 0 568 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_505
timestamp 1554483974
transform 1 0 588 0 1 775
box -3 -3 3 3
use FILL  FILL_597
timestamp 1554483974
transform 1 0 576 0 1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_29
timestamp 1554483974
transform 1 0 584 0 1 770
box -8 -3 104 105
use FILL  FILL_598
timestamp 1554483974
transform 1 0 680 0 1 770
box -8 -3 16 105
use FILL  FILL_599
timestamp 1554483974
transform 1 0 688 0 1 770
box -8 -3 16 105
use FILL  FILL_600
timestamp 1554483974
transform 1 0 696 0 1 770
box -8 -3 16 105
use FILL  FILL_601
timestamp 1554483974
transform 1 0 704 0 1 770
box -8 -3 16 105
use FILL  FILL_602
timestamp 1554483974
transform 1 0 712 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_506
timestamp 1554483974
transform 1 0 732 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_31
timestamp 1554483974
transform 1 0 720 0 1 770
box -8 -3 104 105
use FILL  FILL_604
timestamp 1554483974
transform 1 0 816 0 1 770
box -8 -3 16 105
use FILL  FILL_605
timestamp 1554483974
transform 1 0 824 0 1 770
box -8 -3 16 105
use M3_M2  M3_M2_507
timestamp 1554483974
transform 1 0 844 0 1 775
box -3 -3 3 3
use M3_M2  M3_M2_508
timestamp 1554483974
transform 1 0 868 0 1 775
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_32
timestamp 1554483974
transform 1 0 832 0 1 770
box -8 -3 104 105
use FILL  FILL_606
timestamp 1554483974
transform 1 0 928 0 1 770
box -8 -3 16 105
use FILL  FILL_607
timestamp 1554483974
transform 1 0 936 0 1 770
box -8 -3 16 105
use FILL  FILL_608
timestamp 1554483974
transform 1 0 944 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_11
timestamp 1554483974
transform 1 0 952 0 1 770
box -8 -3 40 105
use FILL  FILL_609
timestamp 1554483974
transform 1 0 984 0 1 770
box -8 -3 16 105
use FILL  FILL_610
timestamp 1554483974
transform 1 0 992 0 1 770
box -8 -3 16 105
use FILL  FILL_624
timestamp 1554483974
transform 1 0 1000 0 1 770
box -8 -3 16 105
use FILL  FILL_626
timestamp 1554483974
transform 1 0 1008 0 1 770
box -8 -3 16 105
use AND2X2  AND2X2_13
timestamp 1554483974
transform 1 0 1016 0 1 770
box -8 -3 40 105
use FILL  FILL_628
timestamp 1554483974
transform 1 0 1048 0 1 770
box -8 -3 16 105
use FILL  FILL_629
timestamp 1554483974
transform 1 0 1056 0 1 770
box -8 -3 16 105
use FILL  FILL_632
timestamp 1554483974
transform 1 0 1064 0 1 770
box -8 -3 16 105
use LATCH  LATCH_10
timestamp 1554483974
transform 1 0 1072 0 1 770
box -8 -3 64 105
use FILL  FILL_634
timestamp 1554483974
transform 1 0 1128 0 1 770
box -8 -3 16 105
use FILL  FILL_640
timestamp 1554483974
transform 1 0 1136 0 1 770
box -8 -3 16 105
use FILL  FILL_642
timestamp 1554483974
transform 1 0 1144 0 1 770
box -8 -3 16 105
use FILL  FILL_644
timestamp 1554483974
transform 1 0 1152 0 1 770
box -8 -3 16 105
use FILL  FILL_645
timestamp 1554483974
transform 1 0 1160 0 1 770
box -8 -3 16 105
use FILL  FILL_646
timestamp 1554483974
transform 1 0 1168 0 1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_27
timestamp 1554483974
transform -1 0 1208 0 1 770
box -8 -3 34 105
use FILL  FILL_647
timestamp 1554483974
transform 1 0 1208 0 1 770
box -8 -3 16 105
use FILL  FILL_649
timestamp 1554483974
transform 1 0 1216 0 1 770
box -8 -3 16 105
use FILL  FILL_651
timestamp 1554483974
transform 1 0 1224 0 1 770
box -8 -3 16 105
use FILL  FILL_653
timestamp 1554483974
transform 1 0 1232 0 1 770
box -8 -3 16 105
use FILL  FILL_654
timestamp 1554483974
transform 1 0 1240 0 1 770
box -8 -3 16 105
use FILL  FILL_655
timestamp 1554483974
transform 1 0 1248 0 1 770
box -8 -3 16 105
use LATCH  LATCH_11
timestamp 1554483974
transform 1 0 1256 0 1 770
box -8 -3 64 105
use FILL  FILL_657
timestamp 1554483974
transform 1 0 1312 0 1 770
box -8 -3 16 105
use FILL  FILL_658
timestamp 1554483974
transform 1 0 1320 0 1 770
box -8 -3 16 105
use FILL  FILL_659
timestamp 1554483974
transform 1 0 1328 0 1 770
box -8 -3 16 105
use LATCH  LATCH_13
timestamp 1554483974
transform 1 0 1336 0 1 770
box -8 -3 64 105
use FILL  FILL_660
timestamp 1554483974
transform 1 0 1392 0 1 770
box -8 -3 16 105
use FILL  FILL_663
timestamp 1554483974
transform 1 0 1400 0 1 770
box -8 -3 16 105
use FILL  FILL_665
timestamp 1554483974
transform 1 0 1408 0 1 770
box -8 -3 16 105
use XOR2X1  XOR2X1_12
timestamp 1554483974
transform 1 0 1416 0 1 770
box -8 -3 64 105
use FILL  FILL_666
timestamp 1554483974
transform 1 0 1472 0 1 770
box -8 -3 16 105
use FILL  FILL_667
timestamp 1554483974
transform 1 0 1480 0 1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_9
timestamp 1554483974
transform 1 0 1488 0 1 770
box -8 -3 40 105
use NOR2X1  NOR2X1_9
timestamp 1554483974
transform 1 0 1520 0 1 770
box -8 -3 32 105
use XOR2X1  XOR2X1_13
timestamp 1554483974
transform 1 0 1544 0 1 770
box -8 -3 64 105
use FILL  FILL_668
timestamp 1554483974
transform 1 0 1600 0 1 770
box -8 -3 16 105
use FILL  FILL_676
timestamp 1554483974
transform 1 0 1608 0 1 770
box -8 -3 16 105
use FILL  FILL_678
timestamp 1554483974
transform 1 0 1616 0 1 770
box -8 -3 16 105
use FILL  FILL_680
timestamp 1554483974
transform 1 0 1624 0 1 770
box -8 -3 16 105
use INVX2  INVX2_43
timestamp 1554483974
transform 1 0 1632 0 1 770
box -9 -3 26 105
use OAI21X1  OAI21X1_29
timestamp 1554483974
transform 1 0 1648 0 1 770
box -8 -3 34 105
use DFFNEGX1  DFFNEGX1_34
timestamp 1554483974
transform 1 0 1680 0 1 770
box -8 -3 104 105
use UART_VIA1  UART_VIA1_17
timestamp 1554483974
transform 1 0 1801 0 1 770
box -10 -3 10 3
use M2_M1  M2_M1_644
timestamp 1554483974
transform 1 0 76 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_645
timestamp 1554483974
transform 1 0 172 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_677
timestamp 1554483974
transform 1 0 84 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_678
timestamp 1554483974
transform 1 0 92 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_679
timestamp 1554483974
transform 1 0 124 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_532
timestamp 1554483974
transform 1 0 172 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_646
timestamp 1554483974
transform 1 0 196 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_680
timestamp 1554483974
transform 1 0 220 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_533
timestamp 1554483974
transform 1 0 268 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_681
timestamp 1554483974
transform 1 0 276 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_682
timestamp 1554483974
transform 1 0 292 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_538
timestamp 1554483974
transform 1 0 276 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_683
timestamp 1554483974
transform 1 0 316 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_684
timestamp 1554483974
transform 1 0 332 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_724
timestamp 1554483974
transform 1 0 324 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_539
timestamp 1554483974
transform 1 0 332 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_737
timestamp 1554483974
transform 1 0 332 0 1 705
box -2 -2 2 2
use M3_M2  M3_M2_540
timestamp 1554483974
transform 1 0 372 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_509
timestamp 1554483974
transform 1 0 404 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_725
timestamp 1554483974
transform 1 0 412 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_726
timestamp 1554483974
transform 1 0 444 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_551
timestamp 1554483974
transform 1 0 444 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_534
timestamp 1554483974
transform 1 0 476 0 1 725
box -3 -3 3 3
use M3_M2  M3_M2_510
timestamp 1554483974
transform 1 0 500 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_520
timestamp 1554483974
transform 1 0 492 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_647
timestamp 1554483974
transform 1 0 500 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_685
timestamp 1554483974
transform 1 0 484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_686
timestamp 1554483974
transform 1 0 492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_687
timestamp 1554483974
transform 1 0 500 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_516
timestamp 1554483974
transform 1 0 532 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_521
timestamp 1554483974
transform 1 0 564 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_688
timestamp 1554483974
transform 1 0 540 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_689
timestamp 1554483974
transform 1 0 556 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_541
timestamp 1554483974
transform 1 0 540 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_727
timestamp 1554483974
transform 1 0 548 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_552
timestamp 1554483974
transform 1 0 548 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_648
timestamp 1554483974
transform 1 0 572 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_553
timestamp 1554483974
transform 1 0 572 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_511
timestamp 1554483974
transform 1 0 676 0 1 765
box -3 -3 3 3
use M3_M2  M3_M2_517
timestamp 1554483974
transform 1 0 588 0 1 755
box -3 -3 3 3
use M3_M2  M3_M2_522
timestamp 1554483974
transform 1 0 636 0 1 745
box -3 -3 3 3
use M3_M2  M3_M2_523
timestamp 1554483974
transform 1 0 692 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_649
timestamp 1554483974
transform 1 0 588 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_526
timestamp 1554483974
transform 1 0 668 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_650
timestamp 1554483974
transform 1 0 676 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_651
timestamp 1554483974
transform 1 0 692 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_527
timestamp 1554483974
transform 1 0 708 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_652
timestamp 1554483974
transform 1 0 716 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_690
timestamp 1554483974
transform 1 0 636 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_691
timestamp 1554483974
transform 1 0 668 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_692
timestamp 1554483974
transform 1 0 684 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_693
timestamp 1554483974
transform 1 0 700 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_542
timestamp 1554483974
transform 1 0 700 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_653
timestamp 1554483974
transform 1 0 796 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_535
timestamp 1554483974
transform 1 0 796 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_654
timestamp 1554483974
transform 1 0 852 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_543
timestamp 1554483974
transform 1 0 852 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_738
timestamp 1554483974
transform 1 0 852 0 1 705
box -2 -2 2 2
use M2_M1  M2_M1_655
timestamp 1554483974
transform 1 0 868 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_656
timestamp 1554483974
transform 1 0 956 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_694
timestamp 1554483974
transform 1 0 892 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_695
timestamp 1554483974
transform 1 0 948 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_544
timestamp 1554483974
transform 1 0 892 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_696
timestamp 1554483974
transform 1 0 972 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_657
timestamp 1554483974
transform 1 0 996 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_528
timestamp 1554483974
transform 1 0 1012 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_697
timestamp 1554483974
transform 1 0 1020 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_561
timestamp 1554483974
transform 1 0 1020 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_698
timestamp 1554483974
transform 1 0 1036 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_545
timestamp 1554483974
transform 1 0 1036 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_658
timestamp 1554483974
transform 1 0 1060 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_546
timestamp 1554483974
transform 1 0 1060 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_529
timestamp 1554483974
transform 1 0 1084 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_699
timestamp 1554483974
transform 1 0 1084 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_554
timestamp 1554483974
transform 1 0 1084 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_700
timestamp 1554483974
transform 1 0 1108 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_536
timestamp 1554483974
transform 1 0 1132 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_728
timestamp 1554483974
transform 1 0 1132 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_524
timestamp 1554483974
transform 1 0 1180 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_659
timestamp 1554483974
transform 1 0 1164 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_660
timestamp 1554483974
transform 1 0 1180 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_701
timestamp 1554483974
transform 1 0 1156 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_702
timestamp 1554483974
transform 1 0 1172 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_703
timestamp 1554483974
transform 1 0 1188 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_525
timestamp 1554483974
transform 1 0 1212 0 1 745
box -3 -3 3 3
use M2_M1  M2_M1_661
timestamp 1554483974
transform 1 0 1204 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_537
timestamp 1554483974
transform 1 0 1204 0 1 725
box -3 -3 3 3
use M2_M1  M2_M1_704
timestamp 1554483974
transform 1 0 1212 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_705
timestamp 1554483974
transform 1 0 1220 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_662
timestamp 1554483974
transform 1 0 1252 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_663
timestamp 1554483974
transform 1 0 1268 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_530
timestamp 1554483974
transform 1 0 1308 0 1 735
box -3 -3 3 3
use M2_M1  M2_M1_664
timestamp 1554483974
transform 1 0 1324 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_665
timestamp 1554483974
transform 1 0 1372 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_706
timestamp 1554483974
transform 1 0 1308 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_729
timestamp 1554483974
transform 1 0 1276 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_555
timestamp 1554483974
transform 1 0 1276 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_707
timestamp 1554483974
transform 1 0 1372 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_708
timestamp 1554483974
transform 1 0 1380 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_730
timestamp 1554483974
transform 1 0 1332 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_562
timestamp 1554483974
transform 1 0 1332 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_512
timestamp 1554483974
transform 1 0 1396 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_666
timestamp 1554483974
transform 1 0 1412 0 1 735
box -2 -2 2 2
use M3_M2  M3_M2_513
timestamp 1554483974
transform 1 0 1460 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_667
timestamp 1554483974
transform 1 0 1444 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_668
timestamp 1554483974
transform 1 0 1460 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_709
timestamp 1554483974
transform 1 0 1420 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_710
timestamp 1554483974
transform 1 0 1436 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_547
timestamp 1554483974
transform 1 0 1420 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_548
timestamp 1554483974
transform 1 0 1444 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_518
timestamp 1554483974
transform 1 0 1492 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_669
timestamp 1554483974
transform 1 0 1492 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_711
timestamp 1554483974
transform 1 0 1468 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_712
timestamp 1554483974
transform 1 0 1484 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_713
timestamp 1554483974
transform 1 0 1492 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_731
timestamp 1554483974
transform 1 0 1460 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_732
timestamp 1554483974
transform 1 0 1468 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_556
timestamp 1554483974
transform 1 0 1468 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_563
timestamp 1554483974
transform 1 0 1460 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_514
timestamp 1554483974
transform 1 0 1524 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_670
timestamp 1554483974
transform 1 0 1524 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_714
timestamp 1554483974
transform 1 0 1516 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_557
timestamp 1554483974
transform 1 0 1516 0 1 705
box -3 -3 3 3
use M3_M2  M3_M2_531
timestamp 1554483974
transform 1 0 1540 0 1 735
box -3 -3 3 3
use M3_M2  M3_M2_519
timestamp 1554483974
transform 1 0 1580 0 1 755
box -3 -3 3 3
use M2_M1  M2_M1_671
timestamp 1554483974
transform 1 0 1564 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_672
timestamp 1554483974
transform 1 0 1580 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_715
timestamp 1554483974
transform 1 0 1556 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_716
timestamp 1554483974
transform 1 0 1572 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_549
timestamp 1554483974
transform 1 0 1540 0 1 715
box -3 -3 3 3
use M3_M2  M3_M2_564
timestamp 1554483974
transform 1 0 1572 0 1 695
box -3 -3 3 3
use M3_M2  M3_M2_515
timestamp 1554483974
transform 1 0 1596 0 1 765
box -3 -3 3 3
use M2_M1  M2_M1_733
timestamp 1554483974
transform 1 0 1596 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_565
timestamp 1554483974
transform 1 0 1596 0 1 695
box -3 -3 3 3
use M2_M1  M2_M1_717
timestamp 1554483974
transform 1 0 1644 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_558
timestamp 1554483974
transform 1 0 1636 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_673
timestamp 1554483974
transform 1 0 1660 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_718
timestamp 1554483974
transform 1 0 1668 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_550
timestamp 1554483974
transform 1 0 1660 0 1 715
box -3 -3 3 3
use M2_M1  M2_M1_734
timestamp 1554483974
transform 1 0 1684 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_735
timestamp 1554483974
transform 1 0 1692 0 1 715
box -2 -2 2 2
use M2_M1  M2_M1_674
timestamp 1554483974
transform 1 0 1700 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_675
timestamp 1554483974
transform 1 0 1724 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_676
timestamp 1554483974
transform 1 0 1732 0 1 735
box -2 -2 2 2
use M2_M1  M2_M1_719
timestamp 1554483974
transform 1 0 1700 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_720
timestamp 1554483974
transform 1 0 1716 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_721
timestamp 1554483974
transform 1 0 1732 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_722
timestamp 1554483974
transform 1 0 1748 0 1 725
box -2 -2 2 2
use M2_M1  M2_M1_723
timestamp 1554483974
transform 1 0 1756 0 1 725
box -2 -2 2 2
use M3_M2  M3_M2_559
timestamp 1554483974
transform 1 0 1692 0 1 705
box -3 -3 3 3
use M2_M1  M2_M1_736
timestamp 1554483974
transform 1 0 1732 0 1 715
box -2 -2 2 2
use M3_M2  M3_M2_560
timestamp 1554483974
transform 1 0 1732 0 1 705
box -3 -3 3 3
use UART_VIA1  UART_VIA1_18
timestamp 1554483974
transform 1 0 24 0 1 670
box -10 -3 10 3
use INVX2  INVX2_34
timestamp 1554483974
transform 1 0 72 0 -1 770
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_27
timestamp 1554483974
transform -1 0 184 0 -1 770
box -8 -3 104 105
use DFFNEGX1  DFFNEGX1_28
timestamp 1554483974
transform 1 0 184 0 -1 770
box -8 -3 104 105
use INVX2  INVX2_35
timestamp 1554483974
transform 1 0 280 0 -1 770
box -9 -3 26 105
use FILL  FILL_562
timestamp 1554483974
transform 1 0 296 0 -1 770
box -8 -3 16 105
use FILL  FILL_563
timestamp 1554483974
transform 1 0 304 0 -1 770
box -8 -3 16 105
use FILL  FILL_564
timestamp 1554483974
transform 1 0 312 0 -1 770
box -8 -3 16 105
use NAND3X1  NAND3X1_7
timestamp 1554483974
transform 1 0 320 0 -1 770
box -8 -3 40 105
use FILL  FILL_565
timestamp 1554483974
transform 1 0 352 0 -1 770
box -8 -3 16 105
use FILL  FILL_566
timestamp 1554483974
transform 1 0 360 0 -1 770
box -8 -3 16 105
use FILL  FILL_567
timestamp 1554483974
transform 1 0 368 0 -1 770
box -8 -3 16 105
use FILL  FILL_569
timestamp 1554483974
transform 1 0 376 0 -1 770
box -8 -3 16 105
use FILL  FILL_571
timestamp 1554483974
transform 1 0 384 0 -1 770
box -8 -3 16 105
use FILL  FILL_573
timestamp 1554483974
transform 1 0 392 0 -1 770
box -8 -3 16 105
use FILL  FILL_577
timestamp 1554483974
transform 1 0 400 0 -1 770
box -8 -3 16 105
use FILL  FILL_578
timestamp 1554483974
transform 1 0 408 0 -1 770
box -8 -3 16 105
use FILL  FILL_579
timestamp 1554483974
transform 1 0 416 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_29
timestamp 1554483974
transform 1 0 424 0 -1 770
box -8 -3 32 105
use FILL  FILL_580
timestamp 1554483974
transform 1 0 448 0 -1 770
box -8 -3 16 105
use FILL  FILL_582
timestamp 1554483974
transform 1 0 456 0 -1 770
box -8 -3 16 105
use FILL  FILL_584
timestamp 1554483974
transform 1 0 464 0 -1 770
box -8 -3 16 105
use FILL  FILL_586
timestamp 1554483974
transform 1 0 472 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_36
timestamp 1554483974
transform 1 0 480 0 -1 770
box -9 -3 26 105
use FILL  FILL_588
timestamp 1554483974
transform 1 0 496 0 -1 770
box -8 -3 16 105
use FILL  FILL_589
timestamp 1554483974
transform 1 0 504 0 -1 770
box -8 -3 16 105
use FILL  FILL_590
timestamp 1554483974
transform 1 0 512 0 -1 770
box -8 -3 16 105
use FILL  FILL_592
timestamp 1554483974
transform 1 0 520 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_31
timestamp 1554483974
transform 1 0 528 0 -1 770
box -8 -3 32 105
use INVX2  INVX2_37
timestamp 1554483974
transform -1 0 568 0 -1 770
box -9 -3 26 105
use FILL  FILL_596
timestamp 1554483974
transform 1 0 568 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_30
timestamp 1554483974
transform 1 0 576 0 -1 770
box -8 -3 104 105
use OAI22X1  OAI22X1_14
timestamp 1554483974
transform -1 0 712 0 -1 770
box -8 -3 46 105
use FILL  FILL_603
timestamp 1554483974
transform 1 0 712 0 -1 770
box -8 -3 16 105
use FILL  FILL_611
timestamp 1554483974
transform 1 0 720 0 -1 770
box -8 -3 16 105
use INVX2  INVX2_38
timestamp 1554483974
transform 1 0 728 0 -1 770
box -9 -3 26 105
use FILL  FILL_612
timestamp 1554483974
transform 1 0 744 0 -1 770
box -8 -3 16 105
use FILL  FILL_613
timestamp 1554483974
transform 1 0 752 0 -1 770
box -8 -3 16 105
use FILL  FILL_614
timestamp 1554483974
transform 1 0 760 0 -1 770
box -8 -3 16 105
use FILL  FILL_615
timestamp 1554483974
transform 1 0 768 0 -1 770
box -8 -3 16 105
use FILL  FILL_616
timestamp 1554483974
transform 1 0 776 0 -1 770
box -8 -3 16 105
use FILL  FILL_617
timestamp 1554483974
transform 1 0 784 0 -1 770
box -8 -3 16 105
use FILL  FILL_618
timestamp 1554483974
transform 1 0 792 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_26
timestamp 1554483974
transform 1 0 800 0 -1 770
box -8 -3 34 105
use FILL  FILL_619
timestamp 1554483974
transform 1 0 832 0 -1 770
box -8 -3 16 105
use FILL  FILL_620
timestamp 1554483974
transform 1 0 840 0 -1 770
box -8 -3 16 105
use FILL  FILL_621
timestamp 1554483974
transform 1 0 848 0 -1 770
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_33
timestamp 1554483974
transform 1 0 856 0 -1 770
box -8 -3 104 105
use FILL  FILL_622
timestamp 1554483974
transform 1 0 952 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_12
timestamp 1554483974
transform 1 0 960 0 -1 770
box -8 -3 40 105
use FILL  FILL_623
timestamp 1554483974
transform 1 0 992 0 -1 770
box -8 -3 16 105
use FILL  FILL_625
timestamp 1554483974
transform 1 0 1000 0 -1 770
box -8 -3 16 105
use FILL  FILL_627
timestamp 1554483974
transform 1 0 1008 0 -1 770
box -8 -3 16 105
use FILL  FILL_630
timestamp 1554483974
transform 1 0 1016 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_14
timestamp 1554483974
transform 1 0 1024 0 -1 770
box -8 -3 40 105
use FILL  FILL_631
timestamp 1554483974
transform 1 0 1056 0 -1 770
box -8 -3 16 105
use FILL  FILL_633
timestamp 1554483974
transform 1 0 1064 0 -1 770
box -8 -3 16 105
use FILL  FILL_635
timestamp 1554483974
transform 1 0 1072 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_32
timestamp 1554483974
transform 1 0 1080 0 -1 770
box -8 -3 32 105
use FILL  FILL_636
timestamp 1554483974
transform 1 0 1104 0 -1 770
box -8 -3 16 105
use FILL  FILL_637
timestamp 1554483974
transform 1 0 1112 0 -1 770
box -8 -3 16 105
use FILL  FILL_638
timestamp 1554483974
transform 1 0 1120 0 -1 770
box -8 -3 16 105
use FILL  FILL_639
timestamp 1554483974
transform 1 0 1128 0 -1 770
box -8 -3 16 105
use FILL  FILL_641
timestamp 1554483974
transform 1 0 1136 0 -1 770
box -8 -3 16 105
use FILL  FILL_643
timestamp 1554483974
transform 1 0 1144 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_5
timestamp 1554483974
transform 1 0 1152 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_39
timestamp 1554483974
transform -1 0 1208 0 -1 770
box -9 -3 26 105
use FILL  FILL_648
timestamp 1554483974
transform 1 0 1208 0 -1 770
box -8 -3 16 105
use FILL  FILL_650
timestamp 1554483974
transform 1 0 1216 0 -1 770
box -8 -3 16 105
use FILL  FILL_652
timestamp 1554483974
transform 1 0 1224 0 -1 770
box -8 -3 16 105
use FILL  FILL_656
timestamp 1554483974
transform 1 0 1232 0 -1 770
box -8 -3 16 105
use M3_M2  M3_M2_566
timestamp 1554483974
transform 1 0 1252 0 1 675
box -3 -3 3 3
use INVX2  INVX2_40
timestamp 1554483974
transform -1 0 1256 0 -1 770
box -9 -3 26 105
use LATCH  LATCH_12
timestamp 1554483974
transform 1 0 1256 0 -1 770
box -8 -3 64 105
use LATCH  LATCH_14
timestamp 1554483974
transform 1 0 1312 0 -1 770
box -8 -3 64 105
use INVX2  INVX2_41
timestamp 1554483974
transform 1 0 1368 0 -1 770
box -9 -3 26 105
use FILL  FILL_661
timestamp 1554483974
transform 1 0 1384 0 -1 770
box -8 -3 16 105
use FILL  FILL_662
timestamp 1554483974
transform 1 0 1392 0 -1 770
box -8 -3 16 105
use FILL  FILL_664
timestamp 1554483974
transform 1 0 1400 0 -1 770
box -8 -3 16 105
use AND2X2  AND2X2_15
timestamp 1554483974
transform 1 0 1408 0 -1 770
box -8 -3 40 105
use NAND2X1  NAND2X1_33
timestamp 1554483974
transform 1 0 1440 0 -1 770
box -8 -3 32 105
use OAI21X1  OAI21X1_28
timestamp 1554483974
transform -1 0 1496 0 -1 770
box -8 -3 34 105
use FILL  FILL_669
timestamp 1554483974
transform 1 0 1496 0 -1 770
box -8 -3 16 105
use FILL  FILL_670
timestamp 1554483974
transform 1 0 1504 0 -1 770
box -8 -3 16 105
use FILL  FILL_671
timestamp 1554483974
transform 1 0 1512 0 -1 770
box -8 -3 16 105
use FILL  FILL_672
timestamp 1554483974
transform 1 0 1520 0 -1 770
box -8 -3 16 105
use FILL  FILL_673
timestamp 1554483974
transform 1 0 1528 0 -1 770
box -8 -3 16 105
use AOI22X1  AOI22X1_6
timestamp 1554483974
transform 1 0 1536 0 -1 770
box -8 -3 46 105
use INVX2  INVX2_42
timestamp 1554483974
transform 1 0 1576 0 -1 770
box -9 -3 26 105
use FILL  FILL_674
timestamp 1554483974
transform 1 0 1592 0 -1 770
box -8 -3 16 105
use FILL  FILL_675
timestamp 1554483974
transform 1 0 1600 0 -1 770
box -8 -3 16 105
use FILL  FILL_677
timestamp 1554483974
transform 1 0 1608 0 -1 770
box -8 -3 16 105
use FILL  FILL_679
timestamp 1554483974
transform 1 0 1616 0 -1 770
box -8 -3 16 105
use FILL  FILL_681
timestamp 1554483974
transform 1 0 1624 0 -1 770
box -8 -3 16 105
use FILL  FILL_682
timestamp 1554483974
transform 1 0 1632 0 -1 770
box -8 -3 16 105
use NAND2X1  NAND2X1_34
timestamp 1554483974
transform -1 0 1664 0 -1 770
box -8 -3 32 105
use NAND2X1  NAND2X1_35
timestamp 1554483974
transform 1 0 1664 0 -1 770
box -8 -3 32 105
use FILL  FILL_683
timestamp 1554483974
transform 1 0 1688 0 -1 770
box -8 -3 16 105
use OAI21X1  OAI21X1_30
timestamp 1554483974
transform -1 0 1728 0 -1 770
box -8 -3 34 105
use OAI21X1  OAI21X1_31
timestamp 1554483974
transform -1 0 1760 0 -1 770
box -8 -3 34 105
use FILL  FILL_684
timestamp 1554483974
transform 1 0 1760 0 -1 770
box -8 -3 16 105
use FILL  FILL_685
timestamp 1554483974
transform 1 0 1768 0 -1 770
box -8 -3 16 105
use UART_VIA1  UART_VIA1_19
timestamp 1554483974
transform 1 0 1825 0 1 670
box -10 -3 10 3
use M3_M2  M3_M2_567
timestamp 1554483974
transform 1 0 92 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_568
timestamp 1554483974
transform 1 0 124 0 1 665
box -3 -3 3 3
use M3_M2  M3_M2_577
timestamp 1554483974
transform 1 0 164 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_589
timestamp 1554483974
transform 1 0 84 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_752
timestamp 1554483974
transform 1 0 108 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_753
timestamp 1554483974
transform 1 0 164 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_754
timestamp 1554483974
transform 1 0 172 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_789
timestamp 1554483974
transform 1 0 84 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_590
timestamp 1554483974
transform 1 0 196 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_755
timestamp 1554483974
transform 1 0 244 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_597
timestamp 1554483974
transform 1 0 244 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_790
timestamp 1554483974
transform 1 0 268 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_571
timestamp 1554483974
transform 1 0 292 0 1 645
box -3 -3 3 3
use M3_M2  M3_M2_578
timestamp 1554483974
transform 1 0 284 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_791
timestamp 1554483974
transform 1 0 284 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_756
timestamp 1554483974
transform 1 0 308 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_572
timestamp 1554483974
transform 1 0 340 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_739
timestamp 1554483974
transform 1 0 340 0 1 635
box -2 -2 2 2
use M3_M2  M3_M2_579
timestamp 1554483974
transform 1 0 324 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_740
timestamp 1554483974
transform 1 0 332 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_580
timestamp 1554483974
transform 1 0 348 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_591
timestamp 1554483974
transform 1 0 332 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_757
timestamp 1554483974
transform 1 0 348 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_598
timestamp 1554483974
transform 1 0 324 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_741
timestamp 1554483974
transform 1 0 372 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_592
timestamp 1554483974
transform 1 0 380 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_742
timestamp 1554483974
transform 1 0 404 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_573
timestamp 1554483974
transform 1 0 428 0 1 645
box -3 -3 3 3
use M2_M1  M2_M1_758
timestamp 1554483974
transform 1 0 420 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_759
timestamp 1554483974
transform 1 0 428 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_792
timestamp 1554483974
transform 1 0 412 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_599
timestamp 1554483974
transform 1 0 420 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_793
timestamp 1554483974
transform 1 0 436 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_600
timestamp 1554483974
transform 1 0 444 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_821
timestamp 1554483974
transform 1 0 444 0 1 595
box -2 -2 2 2
use M3_M2  M3_M2_581
timestamp 1554483974
transform 1 0 476 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_743
timestamp 1554483974
transform 1 0 484 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_760
timestamp 1554483974
transform 1 0 476 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_761
timestamp 1554483974
transform 1 0 484 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_744
timestamp 1554483974
transform 1 0 508 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_794
timestamp 1554483974
transform 1 0 500 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_795
timestamp 1554483974
transform 1 0 524 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_582
timestamp 1554483974
transform 1 0 548 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_745
timestamp 1554483974
transform 1 0 580 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_762
timestamp 1554483974
transform 1 0 564 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_593
timestamp 1554483974
transform 1 0 580 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_796
timestamp 1554483974
transform 1 0 548 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_797
timestamp 1554483974
transform 1 0 556 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_601
timestamp 1554483974
transform 1 0 564 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_583
timestamp 1554483974
transform 1 0 620 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_798
timestamp 1554483974
transform 1 0 620 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_584
timestamp 1554483974
transform 1 0 660 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_763
timestamp 1554483974
transform 1 0 660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_764
timestamp 1554483974
transform 1 0 716 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_765
timestamp 1554483974
transform 1 0 724 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_799
timestamp 1554483974
transform 1 0 636 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_602
timestamp 1554483974
transform 1 0 724 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_607
timestamp 1554483974
transform 1 0 716 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_800
timestamp 1554483974
transform 1 0 748 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_801
timestamp 1554483974
transform 1 0 756 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_608
timestamp 1554483974
transform 1 0 748 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_766
timestamp 1554483974
transform 1 0 812 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_802
timestamp 1554483974
transform 1 0 812 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_609
timestamp 1554483974
transform 1 0 812 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_746
timestamp 1554483974
transform 1 0 828 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_594
timestamp 1554483974
transform 1 0 828 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_767
timestamp 1554483974
transform 1 0 836 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_768
timestamp 1554483974
transform 1 0 844 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_769
timestamp 1554483974
transform 1 0 852 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_603
timestamp 1554483974
transform 1 0 844 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_610
timestamp 1554483974
transform 1 0 836 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_803
timestamp 1554483974
transform 1 0 868 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_604
timestamp 1554483974
transform 1 0 876 0 1 605
box -3 -3 3 3
use M2_M1  M2_M1_747
timestamp 1554483974
transform 1 0 892 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_804
timestamp 1554483974
transform 1 0 932 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_805
timestamp 1554483974
transform 1 0 940 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_574
timestamp 1554483974
transform 1 0 956 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_770
timestamp 1554483974
transform 1 0 956 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_806
timestamp 1554483974
transform 1 0 956 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_611
timestamp 1554483974
transform 1 0 956 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_771
timestamp 1554483974
transform 1 0 972 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_748
timestamp 1554483974
transform 1 0 980 0 1 625
box -2 -2 2 2
use M3_M2  M3_M2_612
timestamp 1554483974
transform 1 0 980 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_772
timestamp 1554483974
transform 1 0 1012 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_605
timestamp 1554483974
transform 1 0 1012 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_595
timestamp 1554483974
transform 1 0 1028 0 1 615
box -3 -3 3 3
use M2_M1  M2_M1_773
timestamp 1554483974
transform 1 0 1044 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_774
timestamp 1554483974
transform 1 0 1052 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_807
timestamp 1554483974
transform 1 0 1028 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_808
timestamp 1554483974
transform 1 0 1036 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_606
timestamp 1554483974
transform 1 0 1052 0 1 605
box -3 -3 3 3
use M3_M2  M3_M2_585
timestamp 1554483974
transform 1 0 1124 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_809
timestamp 1554483974
transform 1 0 1124 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_596
timestamp 1554483974
transform 1 0 1140 0 1 615
box -3 -3 3 3
use M3_M2  M3_M2_586
timestamp 1554483974
transform 1 0 1196 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_775
timestamp 1554483974
transform 1 0 1180 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_776
timestamp 1554483974
transform 1 0 1196 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_810
timestamp 1554483974
transform 1 0 1188 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_613
timestamp 1554483974
transform 1 0 1188 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_777
timestamp 1554483974
transform 1 0 1220 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_575
timestamp 1554483974
transform 1 0 1332 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_778
timestamp 1554483974
transform 1 0 1252 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_779
timestamp 1554483974
transform 1 0 1284 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_811
timestamp 1554483974
transform 1 0 1332 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_614
timestamp 1554483974
transform 1 0 1284 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_576
timestamp 1554483974
transform 1 0 1388 0 1 635
box -3 -3 3 3
use M2_M1  M2_M1_749
timestamp 1554483974
transform 1 0 1404 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_780
timestamp 1554483974
transform 1 0 1388 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_812
timestamp 1554483974
transform 1 0 1380 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_587
timestamp 1554483974
transform 1 0 1428 0 1 625
box -3 -3 3 3
use M3_M2  M3_M2_588
timestamp 1554483974
transform 1 0 1468 0 1 625
box -3 -3 3 3
use M2_M1  M2_M1_781
timestamp 1554483974
transform 1 0 1436 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_782
timestamp 1554483974
transform 1 0 1452 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_783
timestamp 1554483974
transform 1 0 1468 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_813
timestamp 1554483974
transform 1 0 1428 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_814
timestamp 1554483974
transform 1 0 1444 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_815
timestamp 1554483974
transform 1 0 1460 0 1 605
box -2 -2 2 2
use M2_M1  M2_M1_816
timestamp 1554483974
transform 1 0 1476 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_615
timestamp 1554483974
transform 1 0 1444 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_616
timestamp 1554483974
transform 1 0 1468 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_784
timestamp 1554483974
transform 1 0 1492 0 1 615
box -2 -2 2 2
use M3_M2  M3_M2_569
timestamp 1554483974
transform 1 0 1524 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_750
timestamp 1554483974
transform 1 0 1516 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_817
timestamp 1554483974
transform 1 0 1516 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_617
timestamp 1554483974
transform 1 0 1524 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_818
timestamp 1554483974
transform 1 0 1556 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_618
timestamp 1554483974
transform 1 0 1596 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_785
timestamp 1554483974
transform 1 0 1628 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_786
timestamp 1554483974
transform 1 0 1644 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_787
timestamp 1554483974
transform 1 0 1660 0 1 615
box -2 -2 2 2
use M2_M1  M2_M1_819
timestamp 1554483974
transform 1 0 1652 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_619
timestamp 1554483974
transform 1 0 1628 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_570
timestamp 1554483974
transform 1 0 1684 0 1 655
box -3 -3 3 3
use M2_M1  M2_M1_820
timestamp 1554483974
transform 1 0 1684 0 1 605
box -2 -2 2 2
use M3_M2  M3_M2_620
timestamp 1554483974
transform 1 0 1684 0 1 595
box -3 -3 3 3
use M3_M2  M3_M2_621
timestamp 1554483974
transform 1 0 1724 0 1 595
box -3 -3 3 3
use M2_M1  M2_M1_751
timestamp 1554483974
transform 1 0 1748 0 1 625
box -2 -2 2 2
use M2_M1  M2_M1_788
timestamp 1554483974
transform 1 0 1756 0 1 615
box -2 -2 2 2
use UART_VIA1  UART_VIA1_20
timestamp 1554483974
transform 1 0 48 0 1 570
box -10 -3 10 3
use DFFNEGX1  DFFNEGX1_35
timestamp 1554483974
transform 1 0 72 0 1 570
box -8 -3 104 105
use FILL  FILL_686
timestamp 1554483974
transform 1 0 168 0 1 570
box -8 -3 16 105
use FILL  FILL_687
timestamp 1554483974
transform 1 0 176 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_622
timestamp 1554483974
transform 1 0 196 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_36
timestamp 1554483974
transform -1 0 280 0 1 570
box -8 -3 104 105
use FILL  FILL_688
timestamp 1554483974
transform 1 0 280 0 1 570
box -8 -3 16 105
use FILL  FILL_697
timestamp 1554483974
transform 1 0 288 0 1 570
box -8 -3 16 105
use FILL  FILL_699
timestamp 1554483974
transform 1 0 296 0 1 570
box -8 -3 16 105
use FILL  FILL_701
timestamp 1554483974
transform 1 0 304 0 1 570
box -8 -3 16 105
use INVX2  INVX2_44
timestamp 1554483974
transform 1 0 312 0 1 570
box -9 -3 26 105
use NAND3X1  NAND3X1_10
timestamp 1554483974
transform -1 0 360 0 1 570
box -8 -3 40 105
use FILL  FILL_702
timestamp 1554483974
transform 1 0 360 0 1 570
box -8 -3 16 105
use FILL  FILL_704
timestamp 1554483974
transform 1 0 368 0 1 570
box -8 -3 16 105
use FILL  FILL_706
timestamp 1554483974
transform 1 0 376 0 1 570
box -8 -3 16 105
use FILL  FILL_708
timestamp 1554483974
transform 1 0 384 0 1 570
box -8 -3 16 105
use FILL  FILL_710
timestamp 1554483974
transform 1 0 392 0 1 570
box -8 -3 16 105
use FILL  FILL_712
timestamp 1554483974
transform 1 0 400 0 1 570
box -8 -3 16 105
use INVX2  INVX2_46
timestamp 1554483974
transform 1 0 408 0 1 570
box -9 -3 26 105
use NOR2X1  NOR2X1_11
timestamp 1554483974
transform -1 0 448 0 1 570
box -8 -3 32 105
use FILL  FILL_713
timestamp 1554483974
transform 1 0 448 0 1 570
box -8 -3 16 105
use FILL  FILL_714
timestamp 1554483974
transform 1 0 456 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_37
timestamp 1554483974
transform 1 0 464 0 1 570
box -8 -3 32 105
use INVX2  INVX2_48
timestamp 1554483974
transform -1 0 504 0 1 570
box -9 -3 26 105
use FILL  FILL_718
timestamp 1554483974
transform 1 0 504 0 1 570
box -8 -3 16 105
use FILL  FILL_719
timestamp 1554483974
transform 1 0 512 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_32
timestamp 1554483974
transform -1 0 552 0 1 570
box -8 -3 34 105
use M3_M2  M3_M2_623
timestamp 1554483974
transform 1 0 588 0 1 575
box -3 -3 3 3
use OAI21X1  OAI21X1_33
timestamp 1554483974
transform 1 0 552 0 1 570
box -8 -3 34 105
use FILL  FILL_720
timestamp 1554483974
transform 1 0 584 0 1 570
box -8 -3 16 105
use FILL  FILL_722
timestamp 1554483974
transform 1 0 592 0 1 570
box -8 -3 16 105
use FILL  FILL_723
timestamp 1554483974
transform 1 0 600 0 1 570
box -8 -3 16 105
use FILL  FILL_724
timestamp 1554483974
transform 1 0 608 0 1 570
box -8 -3 16 105
use FILL  FILL_725
timestamp 1554483974
transform 1 0 616 0 1 570
box -8 -3 16 105
use M3_M2  M3_M2_624
timestamp 1554483974
transform 1 0 684 0 1 575
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_39
timestamp 1554483974
transform 1 0 624 0 1 570
box -8 -3 104 105
use FILL  FILL_726
timestamp 1554483974
transform 1 0 720 0 1 570
box -8 -3 16 105
use FILL  FILL_727
timestamp 1554483974
transform 1 0 728 0 1 570
box -8 -3 16 105
use INVX2  INVX2_49
timestamp 1554483974
transform -1 0 752 0 1 570
box -9 -3 26 105
use FILL  FILL_728
timestamp 1554483974
transform 1 0 752 0 1 570
box -8 -3 16 105
use FILL  FILL_729
timestamp 1554483974
transform 1 0 760 0 1 570
box -8 -3 16 105
use FILL  FILL_730
timestamp 1554483974
transform 1 0 768 0 1 570
box -8 -3 16 105
use FILL  FILL_731
timestamp 1554483974
transform 1 0 776 0 1 570
box -8 -3 16 105
use FILL  FILL_732
timestamp 1554483974
transform 1 0 784 0 1 570
box -8 -3 16 105
use INVX2  INVX2_50
timestamp 1554483974
transform 1 0 792 0 1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_39
timestamp 1554483974
transform 1 0 808 0 1 570
box -8 -3 32 105
use FILL  FILL_733
timestamp 1554483974
transform 1 0 832 0 1 570
box -8 -3 16 105
use INVX2  INVX2_51
timestamp 1554483974
transform -1 0 856 0 1 570
box -9 -3 26 105
use FILL  FILL_734
timestamp 1554483974
transform 1 0 856 0 1 570
box -8 -3 16 105
use FILL  FILL_735
timestamp 1554483974
transform 1 0 864 0 1 570
box -8 -3 16 105
use FILL  FILL_736
timestamp 1554483974
transform 1 0 872 0 1 570
box -8 -3 16 105
use FILL  FILL_744
timestamp 1554483974
transform 1 0 880 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_40
timestamp 1554483974
transform -1 0 912 0 1 570
box -8 -3 32 105
use FILL  FILL_745
timestamp 1554483974
transform 1 0 912 0 1 570
box -8 -3 16 105
use FILL  FILL_748
timestamp 1554483974
transform 1 0 920 0 1 570
box -8 -3 16 105
use FILL  FILL_750
timestamp 1554483974
transform 1 0 928 0 1 570
box -8 -3 16 105
use INVX2  INVX2_53
timestamp 1554483974
transform 1 0 936 0 1 570
box -9 -3 26 105
use INVX2  INVX2_55
timestamp 1554483974
transform 1 0 952 0 1 570
box -9 -3 26 105
use FILL  FILL_752
timestamp 1554483974
transform 1 0 968 0 1 570
box -8 -3 16 105
use FILL  FILL_756
timestamp 1554483974
transform 1 0 976 0 1 570
box -8 -3 16 105
use FILL  FILL_758
timestamp 1554483974
transform 1 0 984 0 1 570
box -8 -3 16 105
use FILL  FILL_760
timestamp 1554483974
transform 1 0 992 0 1 570
box -8 -3 16 105
use FILL  FILL_762
timestamp 1554483974
transform 1 0 1000 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_41
timestamp 1554483974
transform -1 0 1032 0 1 570
box -8 -3 32 105
use INVX2  INVX2_56
timestamp 1554483974
transform 1 0 1032 0 1 570
box -9 -3 26 105
use FILL  FILL_764
timestamp 1554483974
transform 1 0 1048 0 1 570
box -8 -3 16 105
use FILL  FILL_765
timestamp 1554483974
transform 1 0 1056 0 1 570
box -8 -3 16 105
use FILL  FILL_767
timestamp 1554483974
transform 1 0 1064 0 1 570
box -8 -3 16 105
use FILL  FILL_769
timestamp 1554483974
transform 1 0 1072 0 1 570
box -8 -3 16 105
use FILL  FILL_771
timestamp 1554483974
transform 1 0 1080 0 1 570
box -8 -3 16 105
use FILL  FILL_773
timestamp 1554483974
transform 1 0 1088 0 1 570
box -8 -3 16 105
use FILL  FILL_775
timestamp 1554483974
transform 1 0 1096 0 1 570
box -8 -3 16 105
use FILL  FILL_777
timestamp 1554483974
transform 1 0 1104 0 1 570
box -8 -3 16 105
use INVX2  INVX2_57
timestamp 1554483974
transform -1 0 1128 0 1 570
box -9 -3 26 105
use FILL  FILL_778
timestamp 1554483974
transform 1 0 1128 0 1 570
box -8 -3 16 105
use FILL  FILL_779
timestamp 1554483974
transform 1 0 1136 0 1 570
box -8 -3 16 105
use FILL  FILL_780
timestamp 1554483974
transform 1 0 1144 0 1 570
box -8 -3 16 105
use FILL  FILL_784
timestamp 1554483974
transform 1 0 1152 0 1 570
box -8 -3 16 105
use FILL  FILL_786
timestamp 1554483974
transform 1 0 1160 0 1 570
box -8 -3 16 105
use OAI22X1  OAI22X1_16
timestamp 1554483974
transform -1 0 1208 0 1 570
box -8 -3 46 105
use FILL  FILL_787
timestamp 1554483974
transform 1 0 1208 0 1 570
box -8 -3 16 105
use FILL  FILL_788
timestamp 1554483974
transform 1 0 1216 0 1 570
box -8 -3 16 105
use FILL  FILL_789
timestamp 1554483974
transform 1 0 1224 0 1 570
box -8 -3 16 105
use FILL  FILL_790
timestamp 1554483974
transform 1 0 1232 0 1 570
box -8 -3 16 105
use FILL  FILL_791
timestamp 1554483974
transform 1 0 1240 0 1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_42
timestamp 1554483974
transform -1 0 1344 0 1 570
box -8 -3 104 105
use FILL  FILL_792
timestamp 1554483974
transform 1 0 1344 0 1 570
box -8 -3 16 105
use FILL  FILL_803
timestamp 1554483974
transform 1 0 1352 0 1 570
box -8 -3 16 105
use FILL  FILL_805
timestamp 1554483974
transform 1 0 1360 0 1 570
box -8 -3 16 105
use FILL  FILL_807
timestamp 1554483974
transform 1 0 1368 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_34
timestamp 1554483974
transform 1 0 1376 0 1 570
box -8 -3 34 105
use FILL  FILL_808
timestamp 1554483974
transform 1 0 1408 0 1 570
box -8 -3 16 105
use FILL  FILL_812
timestamp 1554483974
transform 1 0 1416 0 1 570
box -8 -3 16 105
use FILL  FILL_814
timestamp 1554483974
transform 1 0 1424 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_7
timestamp 1554483974
transform 1 0 1432 0 1 570
box -8 -3 46 105
use FILL  FILL_816
timestamp 1554483974
transform 1 0 1472 0 1 570
box -8 -3 16 105
use FILL  FILL_818
timestamp 1554483974
transform 1 0 1480 0 1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_35
timestamp 1554483974
transform 1 0 1488 0 1 570
box -8 -3 34 105
use FILL  FILL_820
timestamp 1554483974
transform 1 0 1520 0 1 570
box -8 -3 16 105
use FILL  FILL_821
timestamp 1554483974
transform 1 0 1528 0 1 570
box -8 -3 16 105
use FILL  FILL_825
timestamp 1554483974
transform 1 0 1536 0 1 570
box -8 -3 16 105
use FILL  FILL_827
timestamp 1554483974
transform 1 0 1544 0 1 570
box -8 -3 16 105
use FILL  FILL_828
timestamp 1554483974
transform 1 0 1552 0 1 570
box -8 -3 16 105
use INVX2  INVX2_60
timestamp 1554483974
transform 1 0 1560 0 1 570
box -9 -3 26 105
use FILL  FILL_829
timestamp 1554483974
transform 1 0 1576 0 1 570
box -8 -3 16 105
use FILL  FILL_830
timestamp 1554483974
transform 1 0 1584 0 1 570
box -8 -3 16 105
use FILL  FILL_833
timestamp 1554483974
transform 1 0 1592 0 1 570
box -8 -3 16 105
use FILL  FILL_835
timestamp 1554483974
transform 1 0 1600 0 1 570
box -8 -3 16 105
use FILL  FILL_837
timestamp 1554483974
transform 1 0 1608 0 1 570
box -8 -3 16 105
use FILL  FILL_839
timestamp 1554483974
transform 1 0 1616 0 1 570
box -8 -3 16 105
use AOI22X1  AOI22X1_8
timestamp 1554483974
transform -1 0 1664 0 1 570
box -8 -3 46 105
use FILL  FILL_840
timestamp 1554483974
transform 1 0 1664 0 1 570
box -8 -3 16 105
use FILL  FILL_845
timestamp 1554483974
transform 1 0 1672 0 1 570
box -8 -3 16 105
use FILL  FILL_847
timestamp 1554483974
transform 1 0 1680 0 1 570
box -8 -3 16 105
use INVX2  INVX2_61
timestamp 1554483974
transform 1 0 1688 0 1 570
box -9 -3 26 105
use FILL  FILL_849
timestamp 1554483974
transform 1 0 1704 0 1 570
box -8 -3 16 105
use FILL  FILL_850
timestamp 1554483974
transform 1 0 1712 0 1 570
box -8 -3 16 105
use FILL  FILL_851
timestamp 1554483974
transform 1 0 1720 0 1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_48
timestamp 1554483974
transform 1 0 1728 0 1 570
box -8 -3 32 105
use FILL  FILL_852
timestamp 1554483974
transform 1 0 1752 0 1 570
box -8 -3 16 105
use FILL  FILL_853
timestamp 1554483974
transform 1 0 1760 0 1 570
box -8 -3 16 105
use FILL  FILL_855
timestamp 1554483974
transform 1 0 1768 0 1 570
box -8 -3 16 105
use UART_VIA1  UART_VIA1_21
timestamp 1554483974
transform 1 0 1801 0 1 570
box -10 -3 10 3
use M2_M1  M2_M1_855
timestamp 1554483974
transform 1 0 76 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_667
timestamp 1554483974
transform 1 0 84 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_630
timestamp 1554483974
transform 1 0 116 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_822
timestamp 1554483974
transform 1 0 116 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_823
timestamp 1554483974
transform 1 0 124 0 1 545
box -2 -2 2 2
use M2_M1  M2_M1_825
timestamp 1554483974
transform 1 0 100 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_826
timestamp 1554483974
transform 1 0 132 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_856
timestamp 1554483974
transform 1 0 116 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_857
timestamp 1554483974
transform 1 0 148 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_827
timestamp 1554483974
transform 1 0 164 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_631
timestamp 1554483974
transform 1 0 204 0 1 555
box -3 -3 3 3
use M2_M1  M2_M1_828
timestamp 1554483974
transform 1 0 252 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_858
timestamp 1554483974
transform 1 0 228 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_654
timestamp 1554483974
transform 1 0 228 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_625
timestamp 1554483974
transform 1 0 268 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_670
timestamp 1554483974
transform 1 0 260 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_859
timestamp 1554483974
transform 1 0 292 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_632
timestamp 1554483974
transform 1 0 340 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_829
timestamp 1554483974
transform 1 0 308 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_830
timestamp 1554483974
transform 1 0 324 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_831
timestamp 1554483974
transform 1 0 340 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_860
timestamp 1554483974
transform 1 0 332 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_861
timestamp 1554483974
transform 1 0 348 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_668
timestamp 1554483974
transform 1 0 308 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_655
timestamp 1554483974
transform 1 0 340 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_671
timestamp 1554483974
transform 1 0 332 0 1 485
box -3 -3 3 3
use M2_M1  M2_M1_832
timestamp 1554483974
transform 1 0 364 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_862
timestamp 1554483974
transform 1 0 356 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_669
timestamp 1554483974
transform 1 0 356 0 1 495
box -3 -3 3 3
use M3_M2  M3_M2_633
timestamp 1554483974
transform 1 0 372 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_833
timestamp 1554483974
transform 1 0 380 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_634
timestamp 1554483974
transform 1 0 420 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_834
timestamp 1554483974
transform 1 0 420 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_635
timestamp 1554483974
transform 1 0 444 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_835
timestamp 1554483974
transform 1 0 436 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_863
timestamp 1554483974
transform 1 0 428 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_836
timestamp 1554483974
transform 1 0 452 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_864
timestamp 1554483974
transform 1 0 444 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_647
timestamp 1554483974
transform 1 0 452 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_663
timestamp 1554483974
transform 1 0 452 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_641
timestamp 1554483974
transform 1 0 476 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_648
timestamp 1554483974
transform 1 0 468 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_626
timestamp 1554483974
transform 1 0 572 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_642
timestamp 1554483974
transform 1 0 508 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_837
timestamp 1554483974
transform 1 0 572 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_865
timestamp 1554483974
transform 1 0 476 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_892
timestamp 1554483974
transform 1 0 468 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_649
timestamp 1554483974
transform 1 0 484 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_866
timestamp 1554483974
transform 1 0 492 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_867
timestamp 1554483974
transform 1 0 524 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_893
timestamp 1554483974
transform 1 0 484 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_664
timestamp 1554483974
transform 1 0 492 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_627
timestamp 1554483974
transform 1 0 596 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_868
timestamp 1554483974
transform 1 0 596 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_628
timestamp 1554483974
transform 1 0 612 0 1 565
box -3 -3 3 3
use M3_M2  M3_M2_629
timestamp 1554483974
transform 1 0 636 0 1 565
box -3 -3 3 3
use M2_M1  M2_M1_869
timestamp 1554483974
transform 1 0 668 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_656
timestamp 1554483974
transform 1 0 668 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_838
timestamp 1554483974
transform 1 0 684 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_870
timestamp 1554483974
transform 1 0 716 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_839
timestamp 1554483974
transform 1 0 860 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_871
timestamp 1554483974
transform 1 0 772 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_872
timestamp 1554483974
transform 1 0 780 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_873
timestamp 1554483974
transform 1 0 836 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_650
timestamp 1554483974
transform 1 0 860 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_874
timestamp 1554483974
transform 1 0 876 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_657
timestamp 1554483974
transform 1 0 876 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_651
timestamp 1554483974
transform 1 0 900 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_875
timestamp 1554483974
transform 1 0 908 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_636
timestamp 1554483974
transform 1 0 948 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_840
timestamp 1554483974
transform 1 0 940 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_876
timestamp 1554483974
transform 1 0 948 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_877
timestamp 1554483974
transform 1 0 956 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_894
timestamp 1554483974
transform 1 0 1012 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_878
timestamp 1554483974
transform 1 0 1036 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_824
timestamp 1554483974
transform 1 0 1052 0 1 545
box -2 -2 2 2
use M3_M2  M3_M2_637
timestamp 1554483974
transform 1 0 1116 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_879
timestamp 1554483974
transform 1 0 1124 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_895
timestamp 1554483974
transform 1 0 1124 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_841
timestamp 1554483974
transform 1 0 1140 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_638
timestamp 1554483974
transform 1 0 1220 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_842
timestamp 1554483974
transform 1 0 1220 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_880
timestamp 1554483974
transform 1 0 1268 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_881
timestamp 1554483974
transform 1 0 1316 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_843
timestamp 1554483974
transform 1 0 1372 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_844
timestamp 1554483974
transform 1 0 1388 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_882
timestamp 1554483974
transform 1 0 1404 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_896
timestamp 1554483974
transform 1 0 1396 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_883
timestamp 1554483974
transform 1 0 1420 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_845
timestamp 1554483974
transform 1 0 1436 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_652
timestamp 1554483974
transform 1 0 1452 0 1 525
box -3 -3 3 3
use M3_M2  M3_M2_658
timestamp 1554483974
transform 1 0 1436 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_846
timestamp 1554483974
transform 1 0 1468 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_884
timestamp 1554483974
transform 1 0 1468 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_665
timestamp 1554483974
transform 1 0 1460 0 1 505
box -3 -3 3 3
use M3_M2  M3_M2_666
timestamp 1554483974
transform 1 0 1476 0 1 505
box -3 -3 3 3
use M2_M1  M2_M1_847
timestamp 1554483974
transform 1 0 1492 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_848
timestamp 1554483974
transform 1 0 1508 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_849
timestamp 1554483974
transform 1 0 1524 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_653
timestamp 1554483974
transform 1 0 1532 0 1 525
box -3 -3 3 3
use M2_M1  M2_M1_897
timestamp 1554483974
transform 1 0 1524 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_898
timestamp 1554483974
transform 1 0 1532 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_643
timestamp 1554483974
transform 1 0 1556 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_885
timestamp 1554483974
transform 1 0 1556 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_850
timestamp 1554483974
transform 1 0 1580 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_644
timestamp 1554483974
transform 1 0 1604 0 1 535
box -3 -3 3 3
use M3_M2  M3_M2_659
timestamp 1554483974
transform 1 0 1604 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_639
timestamp 1554483974
transform 1 0 1620 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_851
timestamp 1554483974
transform 1 0 1620 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_645
timestamp 1554483974
transform 1 0 1644 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_886
timestamp 1554483974
transform 1 0 1628 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_887
timestamp 1554483974
transform 1 0 1636 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_660
timestamp 1554483974
transform 1 0 1636 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_899
timestamp 1554483974
transform 1 0 1652 0 1 515
box -2 -2 2 2
use M2_M1  M2_M1_852
timestamp 1554483974
transform 1 0 1668 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_888
timestamp 1554483974
transform 1 0 1700 0 1 525
box -2 -2 2 2
use M3_M2  M3_M2_661
timestamp 1554483974
transform 1 0 1700 0 1 515
box -3 -3 3 3
use M3_M2  M3_M2_640
timestamp 1554483974
transform 1 0 1756 0 1 545
box -3 -3 3 3
use M2_M1  M2_M1_853
timestamp 1554483974
transform 1 0 1724 0 1 535
box -2 -2 2 2
use M3_M2  M3_M2_646
timestamp 1554483974
transform 1 0 1732 0 1 535
box -3 -3 3 3
use M2_M1  M2_M1_854
timestamp 1554483974
transform 1 0 1756 0 1 535
box -2 -2 2 2
use M2_M1  M2_M1_889
timestamp 1554483974
transform 1 0 1724 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_890
timestamp 1554483974
transform 1 0 1732 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_891
timestamp 1554483974
transform 1 0 1740 0 1 525
box -2 -2 2 2
use M2_M1  M2_M1_900
timestamp 1554483974
transform 1 0 1716 0 1 515
box -2 -2 2 2
use M3_M2  M3_M2_662
timestamp 1554483974
transform 1 0 1732 0 1 515
box -3 -3 3 3
use M2_M1  M2_M1_901
timestamp 1554483974
transform 1 0 1740 0 1 515
box -2 -2 2 2
use UART_VIA1  UART_VIA1_22
timestamp 1554483974
transform 1 0 24 0 1 470
box -10 -3 10 3
use FILL  FILL_689
timestamp 1554483974
transform 1 0 72 0 -1 570
box -8 -3 16 105
use FILL  FILL_690
timestamp 1554483974
transform 1 0 80 0 -1 570
box -8 -3 16 105
use AOI21X1  AOI21X1_1
timestamp 1554483974
transform 1 0 88 0 -1 570
box -7 -3 39 105
use NOR2X1  NOR2X1_10
timestamp 1554483974
transform 1 0 120 0 -1 570
box -8 -3 32 105
use FILL  FILL_691
timestamp 1554483974
transform 1 0 144 0 -1 570
box -8 -3 16 105
use FILL  FILL_692
timestamp 1554483974
transform 1 0 152 0 -1 570
box -8 -3 16 105
use FILL  FILL_693
timestamp 1554483974
transform 1 0 160 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_37
timestamp 1554483974
transform -1 0 264 0 -1 570
box -8 -3 104 105
use FILL  FILL_694
timestamp 1554483974
transform 1 0 264 0 -1 570
box -8 -3 16 105
use FILL  FILL_695
timestamp 1554483974
transform 1 0 272 0 -1 570
box -8 -3 16 105
use FILL  FILL_696
timestamp 1554483974
transform 1 0 280 0 -1 570
box -8 -3 16 105
use FILL  FILL_698
timestamp 1554483974
transform 1 0 288 0 -1 570
box -8 -3 16 105
use FILL  FILL_700
timestamp 1554483974
transform 1 0 296 0 -1 570
box -8 -3 16 105
use M3_M2  M3_M2_672
timestamp 1554483974
transform 1 0 324 0 1 475
box -3 -3 3 3
use M3_M2  M3_M2_673
timestamp 1554483974
transform 1 0 348 0 1 475
box -3 -3 3 3
use OAI22X1  OAI22X1_15
timestamp 1554483974
transform 1 0 304 0 -1 570
box -8 -3 46 105
use INVX2  INVX2_45
timestamp 1554483974
transform -1 0 360 0 -1 570
box -9 -3 26 105
use FILL  FILL_703
timestamp 1554483974
transform 1 0 360 0 -1 570
box -8 -3 16 105
use FILL  FILL_705
timestamp 1554483974
transform 1 0 368 0 -1 570
box -8 -3 16 105
use FILL  FILL_707
timestamp 1554483974
transform 1 0 376 0 -1 570
box -8 -3 16 105
use FILL  FILL_709
timestamp 1554483974
transform 1 0 384 0 -1 570
box -8 -3 16 105
use FILL  FILL_711
timestamp 1554483974
transform 1 0 392 0 -1 570
box -8 -3 16 105
use FILL  FILL_715
timestamp 1554483974
transform 1 0 400 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_47
timestamp 1554483974
transform -1 0 424 0 -1 570
box -9 -3 26 105
use FILL  FILL_716
timestamp 1554483974
transform 1 0 424 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_36
timestamp 1554483974
transform 1 0 432 0 -1 570
box -8 -3 32 105
use FILL  FILL_717
timestamp 1554483974
transform 1 0 456 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_38
timestamp 1554483974
transform 1 0 464 0 -1 570
box -8 -3 32 105
use DFFNEGX1  DFFNEGX1_38
timestamp 1554483974
transform -1 0 584 0 -1 570
box -8 -3 104 105
use FILL  FILL_721
timestamp 1554483974
transform 1 0 584 0 -1 570
box -8 -3 16 105
use FILL  FILL_737
timestamp 1554483974
transform 1 0 592 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_52
timestamp 1554483974
transform -1 0 616 0 -1 570
box -9 -3 26 105
use FILL  FILL_738
timestamp 1554483974
transform 1 0 616 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_0
timestamp 1554483974
transform -1 0 648 0 -1 570
box -5 -3 28 105
use FILL  FILL_739
timestamp 1554483974
transform 1 0 648 0 -1 570
box -8 -3 16 105
use FILL  FILL_740
timestamp 1554483974
transform 1 0 656 0 -1 570
box -8 -3 16 105
use FILL  FILL_741
timestamp 1554483974
transform 1 0 664 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_40
timestamp 1554483974
transform 1 0 672 0 -1 570
box -8 -3 104 105
use FILL  FILL_742
timestamp 1554483974
transform 1 0 768 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_41
timestamp 1554483974
transform -1 0 872 0 -1 570
box -8 -3 104 105
use FILL  FILL_743
timestamp 1554483974
transform 1 0 872 0 -1 570
box -8 -3 16 105
use BUFX2  BUFX2_1
timestamp 1554483974
transform 1 0 880 0 -1 570
box -5 -3 28 105
use FILL  FILL_746
timestamp 1554483974
transform 1 0 904 0 -1 570
box -8 -3 16 105
use FILL  FILL_747
timestamp 1554483974
transform 1 0 912 0 -1 570
box -8 -3 16 105
use FILL  FILL_749
timestamp 1554483974
transform 1 0 920 0 -1 570
box -8 -3 16 105
use FILL  FILL_751
timestamp 1554483974
transform 1 0 928 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_54
timestamp 1554483974
transform 1 0 936 0 -1 570
box -9 -3 26 105
use FILL  FILL_753
timestamp 1554483974
transform 1 0 952 0 -1 570
box -8 -3 16 105
use FILL  FILL_754
timestamp 1554483974
transform 1 0 960 0 -1 570
box -8 -3 16 105
use FILL  FILL_755
timestamp 1554483974
transform 1 0 968 0 -1 570
box -8 -3 16 105
use FILL  FILL_757
timestamp 1554483974
transform 1 0 976 0 -1 570
box -8 -3 16 105
use FILL  FILL_759
timestamp 1554483974
transform 1 0 984 0 -1 570
box -8 -3 16 105
use FILL  FILL_761
timestamp 1554483974
transform 1 0 992 0 -1 570
box -8 -3 16 105
use FILL  FILL_763
timestamp 1554483974
transform 1 0 1000 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_42
timestamp 1554483974
transform -1 0 1032 0 -1 570
box -8 -3 32 105
use NOR2X1  NOR2X1_12
timestamp 1554483974
transform -1 0 1056 0 -1 570
box -8 -3 32 105
use FILL  FILL_766
timestamp 1554483974
transform 1 0 1056 0 -1 570
box -8 -3 16 105
use FILL  FILL_768
timestamp 1554483974
transform 1 0 1064 0 -1 570
box -8 -3 16 105
use FILL  FILL_770
timestamp 1554483974
transform 1 0 1072 0 -1 570
box -8 -3 16 105
use FILL  FILL_772
timestamp 1554483974
transform 1 0 1080 0 -1 570
box -8 -3 16 105
use FILL  FILL_774
timestamp 1554483974
transform 1 0 1088 0 -1 570
box -8 -3 16 105
use FILL  FILL_776
timestamp 1554483974
transform 1 0 1096 0 -1 570
box -8 -3 16 105
use FILL  FILL_781
timestamp 1554483974
transform 1 0 1104 0 -1 570
box -8 -3 16 105
use FILL  FILL_782
timestamp 1554483974
transform 1 0 1112 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_43
timestamp 1554483974
transform -1 0 1144 0 -1 570
box -8 -3 32 105
use FILL  FILL_783
timestamp 1554483974
transform 1 0 1144 0 -1 570
box -8 -3 16 105
use FILL  FILL_785
timestamp 1554483974
transform 1 0 1152 0 -1 570
box -8 -3 16 105
use FILL  FILL_793
timestamp 1554483974
transform 1 0 1160 0 -1 570
box -8 -3 16 105
use FILL  FILL_794
timestamp 1554483974
transform 1 0 1168 0 -1 570
box -8 -3 16 105
use FILL  FILL_795
timestamp 1554483974
transform 1 0 1176 0 -1 570
box -8 -3 16 105
use FILL  FILL_796
timestamp 1554483974
transform 1 0 1184 0 -1 570
box -8 -3 16 105
use FILL  FILL_797
timestamp 1554483974
transform 1 0 1192 0 -1 570
box -8 -3 16 105
use FILL  FILL_798
timestamp 1554483974
transform 1 0 1200 0 -1 570
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_43
timestamp 1554483974
transform 1 0 1208 0 -1 570
box -8 -3 104 105
use INVX2  INVX2_58
timestamp 1554483974
transform 1 0 1304 0 -1 570
box -9 -3 26 105
use FILL  FILL_799
timestamp 1554483974
transform 1 0 1320 0 -1 570
box -8 -3 16 105
use FILL  FILL_800
timestamp 1554483974
transform 1 0 1328 0 -1 570
box -8 -3 16 105
use FILL  FILL_801
timestamp 1554483974
transform 1 0 1336 0 -1 570
box -8 -3 16 105
use FILL  FILL_802
timestamp 1554483974
transform 1 0 1344 0 -1 570
box -8 -3 16 105
use FILL  FILL_804
timestamp 1554483974
transform 1 0 1352 0 -1 570
box -8 -3 16 105
use FILL  FILL_806
timestamp 1554483974
transform 1 0 1360 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_44
timestamp 1554483974
transform 1 0 1368 0 -1 570
box -8 -3 32 105
use FILL  FILL_809
timestamp 1554483974
transform 1 0 1392 0 -1 570
box -8 -3 16 105
use FILL  FILL_810
timestamp 1554483974
transform 1 0 1400 0 -1 570
box -8 -3 16 105
use FILL  FILL_811
timestamp 1554483974
transform 1 0 1408 0 -1 570
box -8 -3 16 105
use FILL  FILL_813
timestamp 1554483974
transform 1 0 1416 0 -1 570
box -8 -3 16 105
use FILL  FILL_815
timestamp 1554483974
transform 1 0 1424 0 -1 570
box -8 -3 16 105
use INVX2  INVX2_59
timestamp 1554483974
transform 1 0 1432 0 -1 570
box -9 -3 26 105
use NAND2X1  NAND2X1_45
timestamp 1554483974
transform -1 0 1472 0 -1 570
box -8 -3 32 105
use FILL  FILL_817
timestamp 1554483974
transform 1 0 1472 0 -1 570
box -8 -3 16 105
use FILL  FILL_819
timestamp 1554483974
transform 1 0 1480 0 -1 570
box -8 -3 16 105
use FILL  FILL_822
timestamp 1554483974
transform 1 0 1488 0 -1 570
box -8 -3 16 105
use FILL  FILL_823
timestamp 1554483974
transform 1 0 1496 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_46
timestamp 1554483974
transform 1 0 1504 0 -1 570
box -8 -3 32 105
use FILL  FILL_824
timestamp 1554483974
transform 1 0 1528 0 -1 570
box -8 -3 16 105
use FILL  FILL_826
timestamp 1554483974
transform 1 0 1536 0 -1 570
box -8 -3 16 105
use FILL  FILL_831
timestamp 1554483974
transform 1 0 1544 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_36
timestamp 1554483974
transform -1 0 1584 0 -1 570
box -8 -3 34 105
use FILL  FILL_832
timestamp 1554483974
transform 1 0 1584 0 -1 570
box -8 -3 16 105
use FILL  FILL_834
timestamp 1554483974
transform 1 0 1592 0 -1 570
box -8 -3 16 105
use FILL  FILL_836
timestamp 1554483974
transform 1 0 1600 0 -1 570
box -8 -3 16 105
use FILL  FILL_838
timestamp 1554483974
transform 1 0 1608 0 -1 570
box -8 -3 16 105
use FILL  FILL_841
timestamp 1554483974
transform 1 0 1616 0 -1 570
box -8 -3 16 105
use FILL  FILL_842
timestamp 1554483974
transform 1 0 1624 0 -1 570
box -8 -3 16 105
use NAND2X1  NAND2X1_47
timestamp 1554483974
transform 1 0 1632 0 -1 570
box -8 -3 32 105
use FILL  FILL_843
timestamp 1554483974
transform 1 0 1656 0 -1 570
box -8 -3 16 105
use FILL  FILL_844
timestamp 1554483974
transform 1 0 1664 0 -1 570
box -8 -3 16 105
use FILL  FILL_846
timestamp 1554483974
transform 1 0 1672 0 -1 570
box -8 -3 16 105
use FILL  FILL_848
timestamp 1554483974
transform 1 0 1680 0 -1 570
box -8 -3 16 105
use OAI21X1  OAI21X1_37
timestamp 1554483974
transform 1 0 1688 0 -1 570
box -8 -3 34 105
use NAND2X1  NAND2X1_49
timestamp 1554483974
transform 1 0 1720 0 -1 570
box -8 -3 32 105
use M3_M2  M3_M2_674
timestamp 1554483974
transform 1 0 1756 0 1 475
box -3 -3 3 3
use INVX2  INVX2_62
timestamp 1554483974
transform -1 0 1760 0 -1 570
box -9 -3 26 105
use M3_M2  M3_M2_675
timestamp 1554483974
transform 1 0 1772 0 1 475
box -3 -3 3 3
use FILL  FILL_854
timestamp 1554483974
transform 1 0 1760 0 -1 570
box -8 -3 16 105
use FILL  FILL_856
timestamp 1554483974
transform 1 0 1768 0 -1 570
box -8 -3 16 105
use UART_VIA1  UART_VIA1_23
timestamp 1554483974
transform 1 0 1825 0 1 470
box -10 -3 10 3
use M2_M1  M2_M1_905
timestamp 1554483974
transform 1 0 100 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_902
timestamp 1554483974
transform 1 0 132 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_906
timestamp 1554483974
transform 1 0 132 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_913
timestamp 1554483974
transform 1 0 124 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_699
timestamp 1554483974
transform 1 0 132 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_907
timestamp 1554483974
transform 1 0 148 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_914
timestamp 1554483974
transform 1 0 180 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_709
timestamp 1554483974
transform 1 0 180 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_679
timestamp 1554483974
transform 1 0 204 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_949
timestamp 1554483974
transform 1 0 188 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_710
timestamp 1554483974
transform 1 0 212 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_981
timestamp 1554483974
transform 1 0 204 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_915
timestamp 1554483974
transform 1 0 220 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_700
timestamp 1554483974
transform 1 0 236 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_950
timestamp 1554483974
transform 1 0 236 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_916
timestamp 1554483974
transform 1 0 252 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_718
timestamp 1554483974
transform 1 0 252 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_701
timestamp 1554483974
transform 1 0 268 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_951
timestamp 1554483974
transform 1 0 308 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_917
timestamp 1554483974
transform 1 0 324 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_918
timestamp 1554483974
transform 1 0 348 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_680
timestamp 1554483974
transform 1 0 364 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_919
timestamp 1554483974
transform 1 0 364 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_952
timestamp 1554483974
transform 1 0 340 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_953
timestamp 1554483974
transform 1 0 356 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_719
timestamp 1554483974
transform 1 0 348 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_954
timestamp 1554483974
transform 1 0 372 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_920
timestamp 1554483974
transform 1 0 396 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_921
timestamp 1554483974
transform 1 0 444 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_955
timestamp 1554483974
transform 1 0 420 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_956
timestamp 1554483974
transform 1 0 428 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_720
timestamp 1554483974
transform 1 0 420 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_982
timestamp 1554483974
transform 1 0 428 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_728
timestamp 1554483974
transform 1 0 428 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_729
timestamp 1554483974
transform 1 0 444 0 1 385
box -3 -3 3 3
use M3_M2  M3_M2_688
timestamp 1554483974
transform 1 0 468 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_689
timestamp 1554483974
transform 1 0 508 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_922
timestamp 1554483974
transform 1 0 468 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_923
timestamp 1554483974
transform 1 0 476 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_924
timestamp 1554483974
transform 1 0 508 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_957
timestamp 1554483974
transform 1 0 556 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_730
timestamp 1554483974
transform 1 0 476 0 1 385
box -3 -3 3 3
use M2_M1  M2_M1_925
timestamp 1554483974
transform 1 0 620 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_958
timestamp 1554483974
transform 1 0 588 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_721
timestamp 1554483974
transform 1 0 668 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_681
timestamp 1554483974
transform 1 0 700 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_926
timestamp 1554483974
transform 1 0 700 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_927
timestamp 1554483974
transform 1 0 708 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_676
timestamp 1554483974
transform 1 0 772 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_928
timestamp 1554483974
transform 1 0 740 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_929
timestamp 1554483974
transform 1 0 796 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_702
timestamp 1554483974
transform 1 0 820 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_930
timestamp 1554483974
transform 1 0 836 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_931
timestamp 1554483974
transform 1 0 852 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_959
timestamp 1554483974
transform 1 0 724 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_711
timestamp 1554483974
transform 1 0 732 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_712
timestamp 1554483974
transform 1 0 780 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_960
timestamp 1554483974
transform 1 0 820 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_722
timestamp 1554483974
transform 1 0 724 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_983
timestamp 1554483974
transform 1 0 732 0 1 395
box -2 -2 2 2
use M3_M2  M3_M2_723
timestamp 1554483974
transform 1 0 756 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_724
timestamp 1554483974
transform 1 0 796 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_703
timestamp 1554483974
transform 1 0 860 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_713
timestamp 1554483974
transform 1 0 852 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_714
timestamp 1554483974
transform 1 0 892 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_682
timestamp 1554483974
transform 1 0 908 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_961
timestamp 1554483974
transform 1 0 900 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_962
timestamp 1554483974
transform 1 0 908 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_690
timestamp 1554483974
transform 1 0 916 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_932
timestamp 1554483974
transform 1 0 916 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_933
timestamp 1554483974
transform 1 0 924 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_691
timestamp 1554483974
transform 1 0 940 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_715
timestamp 1554483974
transform 1 0 932 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_725
timestamp 1554483974
transform 1 0 932 0 1 395
box -3 -3 3 3
use M2_M1  M2_M1_963
timestamp 1554483974
transform 1 0 948 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_934
timestamp 1554483974
transform 1 0 956 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_964
timestamp 1554483974
transform 1 0 964 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_677
timestamp 1554483974
transform 1 0 980 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_903
timestamp 1554483974
transform 1 0 980 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_908
timestamp 1554483974
transform 1 0 980 0 1 425
box -2 -2 2 2
use M3_M2  M3_M2_683
timestamp 1554483974
transform 1 0 1020 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_692
timestamp 1554483974
transform 1 0 1012 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_909
timestamp 1554483974
transform 1 0 1028 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_935
timestamp 1554483974
transform 1 0 1012 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_936
timestamp 1554483974
transform 1 0 1036 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_693
timestamp 1554483974
transform 1 0 1076 0 1 425
box -3 -3 3 3
use M3_M2  M3_M2_704
timestamp 1554483974
transform 1 0 1068 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_678
timestamp 1554483974
transform 1 0 1100 0 1 445
box -3 -3 3 3
use M2_M1  M2_M1_904
timestamp 1554483974
transform 1 0 1100 0 1 435
box -2 -2 2 2
use M2_M1  M2_M1_910
timestamp 1554483974
transform 1 0 1100 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_965
timestamp 1554483974
transform 1 0 1092 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_694
timestamp 1554483974
transform 1 0 1124 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_911
timestamp 1554483974
transform 1 0 1140 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_937
timestamp 1554483974
transform 1 0 1124 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_705
timestamp 1554483974
transform 1 0 1148 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_912
timestamp 1554483974
transform 1 0 1164 0 1 425
box -2 -2 2 2
use M2_M1  M2_M1_938
timestamp 1554483974
transform 1 0 1156 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_966
timestamp 1554483974
transform 1 0 1148 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_706
timestamp 1554483974
transform 1 0 1164 0 1 415
box -3 -3 3 3
use M3_M2  M3_M2_684
timestamp 1554483974
transform 1 0 1252 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_939
timestamp 1554483974
transform 1 0 1252 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_967
timestamp 1554483974
transform 1 0 1244 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_968
timestamp 1554483974
transform 1 0 1252 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_685
timestamp 1554483974
transform 1 0 1284 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_695
timestamp 1554483974
transform 1 0 1268 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_940
timestamp 1554483974
transform 1 0 1268 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_941
timestamp 1554483974
transform 1 0 1284 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_969
timestamp 1554483974
transform 1 0 1276 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_970
timestamp 1554483974
transform 1 0 1316 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_696
timestamp 1554483974
transform 1 0 1332 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_971
timestamp 1554483974
transform 1 0 1332 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_972
timestamp 1554483974
transform 1 0 1428 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_973
timestamp 1554483974
transform 1 0 1452 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_974
timestamp 1554483974
transform 1 0 1460 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_707
timestamp 1554483974
transform 1 0 1484 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_984
timestamp 1554483974
transform 1 0 1484 0 1 395
box -2 -2 2 2
use M2_M1  M2_M1_942
timestamp 1554483974
transform 1 0 1500 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_943
timestamp 1554483974
transform 1 0 1508 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_708
timestamp 1554483974
transform 1 0 1524 0 1 415
box -3 -3 3 3
use M2_M1  M2_M1_975
timestamp 1554483974
transform 1 0 1524 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_716
timestamp 1554483974
transform 1 0 1532 0 1 405
box -3 -3 3 3
use M3_M2  M3_M2_686
timestamp 1554483974
transform 1 0 1596 0 1 435
box -3 -3 3 3
use M2_M1  M2_M1_944
timestamp 1554483974
transform 1 0 1612 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_945
timestamp 1554483974
transform 1 0 1644 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_976
timestamp 1554483974
transform 1 0 1604 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_717
timestamp 1554483974
transform 1 0 1612 0 1 405
box -3 -3 3 3
use M2_M1  M2_M1_977
timestamp 1554483974
transform 1 0 1620 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_978
timestamp 1554483974
transform 1 0 1636 0 1 405
box -2 -2 2 2
use M2_M1  M2_M1_979
timestamp 1554483974
transform 1 0 1644 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_726
timestamp 1554483974
transform 1 0 1620 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_727
timestamp 1554483974
transform 1 0 1644 0 1 395
box -3 -3 3 3
use M3_M2  M3_M2_697
timestamp 1554483974
transform 1 0 1676 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_946
timestamp 1554483974
transform 1 0 1676 0 1 415
box -2 -2 2 2
use M3_M2  M3_M2_687
timestamp 1554483974
transform 1 0 1780 0 1 435
box -3 -3 3 3
use M3_M2  M3_M2_698
timestamp 1554483974
transform 1 0 1716 0 1 425
box -3 -3 3 3
use M2_M1  M2_M1_947
timestamp 1554483974
transform 1 0 1724 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_948
timestamp 1554483974
transform 1 0 1772 0 1 415
box -2 -2 2 2
use M2_M1  M2_M1_980
timestamp 1554483974
transform 1 0 1692 0 1 405
box -2 -2 2 2
use M3_M2  M3_M2_731
timestamp 1554483974
transform 1 0 1772 0 1 385
box -3 -3 3 3
use UART_VIA1  UART_VIA1_24
timestamp 1554483974
transform 1 0 48 0 1 370
box -10 -3 10 3
use FILL  FILL_857
timestamp 1554483974
transform 1 0 72 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_732
timestamp 1554483974
transform 1 0 92 0 1 375
box -3 -3 3 3
use FILL  FILL_859
timestamp 1554483974
transform 1 0 80 0 1 370
box -8 -3 16 105
use FILL  FILL_861
timestamp 1554483974
transform 1 0 88 0 1 370
box -8 -3 16 105
use FILL  FILL_863
timestamp 1554483974
transform 1 0 96 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_11
timestamp 1554483974
transform -1 0 136 0 1 370
box -8 -3 40 105
use FILL  FILL_864
timestamp 1554483974
transform 1 0 136 0 1 370
box -8 -3 16 105
use FILL  FILL_871
timestamp 1554483974
transform 1 0 144 0 1 370
box -8 -3 16 105
use M3_M2  M3_M2_733
timestamp 1554483974
transform 1 0 164 0 1 375
box -3 -3 3 3
use FILL  FILL_873
timestamp 1554483974
transform 1 0 152 0 1 370
box -8 -3 16 105
use FILL  FILL_875
timestamp 1554483974
transform 1 0 160 0 1 370
box -8 -3 16 105
use FILL  FILL_876
timestamp 1554483974
transform 1 0 168 0 1 370
box -8 -3 16 105
use AOI21X1  AOI21X1_2
timestamp 1554483974
transform 1 0 176 0 1 370
box -7 -3 39 105
use FILL  FILL_877
timestamp 1554483974
transform 1 0 208 0 1 370
box -8 -3 16 105
use FILL  FILL_881
timestamp 1554483974
transform 1 0 216 0 1 370
box -8 -3 16 105
use FILL  FILL_883
timestamp 1554483974
transform 1 0 224 0 1 370
box -8 -3 16 105
use FILL  FILL_885
timestamp 1554483974
transform 1 0 232 0 1 370
box -8 -3 16 105
use INVX2  INVX2_63
timestamp 1554483974
transform 1 0 240 0 1 370
box -9 -3 26 105
use FILL  FILL_886
timestamp 1554483974
transform 1 0 256 0 1 370
box -8 -3 16 105
use FILL  FILL_887
timestamp 1554483974
transform 1 0 264 0 1 370
box -8 -3 16 105
use FILL  FILL_888
timestamp 1554483974
transform 1 0 272 0 1 370
box -8 -3 16 105
use FILL  FILL_891
timestamp 1554483974
transform 1 0 280 0 1 370
box -8 -3 16 105
use FILL  FILL_893
timestamp 1554483974
transform 1 0 288 0 1 370
box -8 -3 16 105
use FILL  FILL_895
timestamp 1554483974
transform 1 0 296 0 1 370
box -8 -3 16 105
use FILL  FILL_897
timestamp 1554483974
transform 1 0 304 0 1 370
box -8 -3 16 105
use FILL  FILL_899
timestamp 1554483974
transform 1 0 312 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_17
timestamp 1554483974
transform 1 0 320 0 1 370
box -8 -3 46 105
use FILL  FILL_901
timestamp 1554483974
transform 1 0 360 0 1 370
box -8 -3 16 105
use FILL  FILL_903
timestamp 1554483974
transform 1 0 368 0 1 370
box -8 -3 16 105
use FILL  FILL_905
timestamp 1554483974
transform 1 0 376 0 1 370
box -8 -3 16 105
use FILL  FILL_907
timestamp 1554483974
transform 1 0 384 0 1 370
box -8 -3 16 105
use FILL  FILL_909
timestamp 1554483974
transform 1 0 392 0 1 370
box -8 -3 16 105
use OR2X1  OR2X1_2
timestamp 1554483974
transform -1 0 432 0 1 370
box -8 -3 40 105
use AND2X2  AND2X2_16
timestamp 1554483974
transform 1 0 432 0 1 370
box -8 -3 40 105
use FILL  FILL_910
timestamp 1554483974
transform 1 0 464 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_44
timestamp 1554483974
transform -1 0 568 0 1 370
box -8 -3 104 105
use FILL  FILL_911
timestamp 1554483974
transform 1 0 568 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_45
timestamp 1554483974
transform 1 0 576 0 1 370
box -8 -3 104 105
use FILL  FILL_912
timestamp 1554483974
transform 1 0 672 0 1 370
box -8 -3 16 105
use FILL  FILL_922
timestamp 1554483974
transform 1 0 680 0 1 370
box -8 -3 16 105
use FILL  FILL_924
timestamp 1554483974
transform 1 0 688 0 1 370
box -8 -3 16 105
use FILL  FILL_925
timestamp 1554483974
transform 1 0 696 0 1 370
box -8 -3 16 105
use OR2X1  OR2X1_3
timestamp 1554483974
transform -1 0 736 0 1 370
box -8 -3 40 105
use DFFNEGX1  DFFNEGX1_48
timestamp 1554483974
transform -1 0 832 0 1 370
box -8 -3 104 105
use AND2X2  AND2X2_17
timestamp 1554483974
transform -1 0 864 0 1 370
box -8 -3 40 105
use FILL  FILL_926
timestamp 1554483974
transform 1 0 864 0 1 370
box -8 -3 16 105
use FILL  FILL_942
timestamp 1554483974
transform 1 0 872 0 1 370
box -8 -3 16 105
use FILL  FILL_944
timestamp 1554483974
transform 1 0 880 0 1 370
box -8 -3 16 105
use FILL  FILL_946
timestamp 1554483974
transform 1 0 888 0 1 370
box -8 -3 16 105
use FILL  FILL_948
timestamp 1554483974
transform 1 0 896 0 1 370
box -8 -3 16 105
use INVX2  INVX2_64
timestamp 1554483974
transform 1 0 904 0 1 370
box -9 -3 26 105
use INVX2  INVX2_65
timestamp 1554483974
transform -1 0 936 0 1 370
box -9 -3 26 105
use FILL  FILL_950
timestamp 1554483974
transform 1 0 936 0 1 370
box -8 -3 16 105
use FILL  FILL_951
timestamp 1554483974
transform 1 0 944 0 1 370
box -8 -3 16 105
use FILL  FILL_952
timestamp 1554483974
transform 1 0 952 0 1 370
box -8 -3 16 105
use INVX2  INVX2_66
timestamp 1554483974
transform 1 0 960 0 1 370
box -9 -3 26 105
use FILL  FILL_955
timestamp 1554483974
transform 1 0 976 0 1 370
box -8 -3 16 105
use FILL  FILL_959
timestamp 1554483974
transform 1 0 984 0 1 370
box -8 -3 16 105
use FILL  FILL_961
timestamp 1554483974
transform 1 0 992 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_15
timestamp 1554483974
transform 1 0 1000 0 1 370
box -8 -3 40 105
use FILL  FILL_963
timestamp 1554483974
transform 1 0 1032 0 1 370
box -8 -3 16 105
use FILL  FILL_964
timestamp 1554483974
transform 1 0 1040 0 1 370
box -8 -3 16 105
use FILL  FILL_965
timestamp 1554483974
transform 1 0 1048 0 1 370
box -8 -3 16 105
use FILL  FILL_969
timestamp 1554483974
transform 1 0 1056 0 1 370
box -8 -3 16 105
use FILL  FILL_971
timestamp 1554483974
transform 1 0 1064 0 1 370
box -8 -3 16 105
use FILL  FILL_973
timestamp 1554483974
transform 1 0 1072 0 1 370
box -8 -3 16 105
use INVX2  INVX2_67
timestamp 1554483974
transform -1 0 1096 0 1 370
box -9 -3 26 105
use FILL  FILL_974
timestamp 1554483974
transform 1 0 1096 0 1 370
box -8 -3 16 105
use FILL  FILL_975
timestamp 1554483974
transform 1 0 1104 0 1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_18
timestamp 1554483974
transform 1 0 1112 0 1 370
box -8 -3 40 105
use INVX2  INVX2_68
timestamp 1554483974
transform 1 0 1144 0 1 370
box -9 -3 26 105
use FILL  FILL_977
timestamp 1554483974
transform 1 0 1160 0 1 370
box -8 -3 16 105
use FILL  FILL_978
timestamp 1554483974
transform 1 0 1168 0 1 370
box -8 -3 16 105
use FILL  FILL_979
timestamp 1554483974
transform 1 0 1176 0 1 370
box -8 -3 16 105
use FILL  FILL_980
timestamp 1554483974
transform 1 0 1184 0 1 370
box -8 -3 16 105
use FILL  FILL_981
timestamp 1554483974
transform 1 0 1192 0 1 370
box -8 -3 16 105
use FILL  FILL_982
timestamp 1554483974
transform 1 0 1200 0 1 370
box -8 -3 16 105
use FILL  FILL_983
timestamp 1554483974
transform 1 0 1208 0 1 370
box -8 -3 16 105
use FILL  FILL_984
timestamp 1554483974
transform 1 0 1216 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_50
timestamp 1554483974
transform -1 0 1248 0 1 370
box -8 -3 32 105
use FILL  FILL_985
timestamp 1554483974
transform 1 0 1248 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_20
timestamp 1554483974
transform -1 0 1296 0 1 370
box -8 -3 46 105
use FILL  FILL_986
timestamp 1554483974
transform 1 0 1296 0 1 370
box -8 -3 16 105
use FILL  FILL_987
timestamp 1554483974
transform 1 0 1304 0 1 370
box -8 -3 16 105
use FILL  FILL_988
timestamp 1554483974
transform 1 0 1312 0 1 370
box -8 -3 16 105
use FILL  FILL_1003
timestamp 1554483974
transform 1 0 1320 0 1 370
box -8 -3 16 105
use FILL  FILL_1005
timestamp 1554483974
transform 1 0 1328 0 1 370
box -8 -3 16 105
use OAI21X1  OAI21X1_39
timestamp 1554483974
transform -1 0 1368 0 1 370
box -8 -3 34 105
use FILL  FILL_1006
timestamp 1554483974
transform 1 0 1368 0 1 370
box -8 -3 16 105
use FILL  FILL_1007
timestamp 1554483974
transform 1 0 1376 0 1 370
box -8 -3 16 105
use FILL  FILL_1012
timestamp 1554483974
transform 1 0 1384 0 1 370
box -8 -3 16 105
use FILL  FILL_1014
timestamp 1554483974
transform 1 0 1392 0 1 370
box -8 -3 16 105
use FILL  FILL_1016
timestamp 1554483974
transform 1 0 1400 0 1 370
box -8 -3 16 105
use FILL  FILL_1018
timestamp 1554483974
transform 1 0 1408 0 1 370
box -8 -3 16 105
use FILL  FILL_1020
timestamp 1554483974
transform 1 0 1416 0 1 370
box -8 -3 16 105
use FILL  FILL_1021
timestamp 1554483974
transform 1 0 1424 0 1 370
box -8 -3 16 105
use OR2X1  OR2X1_4
timestamp 1554483974
transform -1 0 1464 0 1 370
box -8 -3 40 105
use FILL  FILL_1022
timestamp 1554483974
transform 1 0 1464 0 1 370
box -8 -3 16 105
use FILL  FILL_1025
timestamp 1554483974
transform 1 0 1472 0 1 370
box -8 -3 16 105
use FILL  FILL_1027
timestamp 1554483974
transform 1 0 1480 0 1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_54
timestamp 1554483974
transform 1 0 1488 0 1 370
box -8 -3 32 105
use INVX2  INVX2_71
timestamp 1554483974
transform -1 0 1528 0 1 370
box -9 -3 26 105
use FILL  FILL_1029
timestamp 1554483974
transform 1 0 1528 0 1 370
box -8 -3 16 105
use FILL  FILL_1032
timestamp 1554483974
transform 1 0 1536 0 1 370
box -8 -3 16 105
use FILL  FILL_1034
timestamp 1554483974
transform 1 0 1544 0 1 370
box -8 -3 16 105
use FILL  FILL_1036
timestamp 1554483974
transform 1 0 1552 0 1 370
box -8 -3 16 105
use FILL  FILL_1038
timestamp 1554483974
transform 1 0 1560 0 1 370
box -8 -3 16 105
use FILL  FILL_1039
timestamp 1554483974
transform 1 0 1568 0 1 370
box -8 -3 16 105
use FILL  FILL_1040
timestamp 1554483974
transform 1 0 1576 0 1 370
box -8 -3 16 105
use FILL  FILL_1041
timestamp 1554483974
transform 1 0 1584 0 1 370
box -8 -3 16 105
use FILL  FILL_1042
timestamp 1554483974
transform 1 0 1592 0 1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_21
timestamp 1554483974
transform -1 0 1640 0 1 370
box -8 -3 46 105
use INVX2  INVX2_72
timestamp 1554483974
transform 1 0 1640 0 1 370
box -9 -3 26 105
use FILL  FILL_1043
timestamp 1554483974
transform 1 0 1656 0 1 370
box -8 -3 16 105
use FILL  FILL_1044
timestamp 1554483974
transform 1 0 1664 0 1 370
box -8 -3 16 105
use FILL  FILL_1045
timestamp 1554483974
transform 1 0 1672 0 1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_49
timestamp 1554483974
transform 1 0 1680 0 1 370
box -8 -3 104 105
use UART_VIA1  UART_VIA1_25
timestamp 1554483974
transform 1 0 1801 0 1 370
box -10 -3 10 3
use M2_M1  M2_M1_1055
timestamp 1554483974
transform 1 0 92 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_760
timestamp 1554483974
transform 1 0 108 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1041
timestamp 1554483974
transform 1 0 124 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1056
timestamp 1554483974
transform 1 0 132 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_761
timestamp 1554483974
transform 1 0 164 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1015
timestamp 1554483974
transform 1 0 172 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1042
timestamp 1554483974
transform 1 0 172 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1043
timestamp 1554483974
transform 1 0 188 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_771
timestamp 1554483974
transform 1 0 172 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_1044
timestamp 1554483974
transform 1 0 212 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_762
timestamp 1554483974
transform 1 0 252 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1016
timestamp 1554483974
transform 1 0 260 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1045
timestamp 1554483974
transform 1 0 268 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1057
timestamp 1554483974
transform 1 0 268 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1017
timestamp 1554483974
transform 1 0 292 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_988
timestamp 1554483974
transform 1 0 308 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_989
timestamp 1554483974
transform 1 0 340 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_990
timestamp 1554483974
transform 1 0 356 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1018
timestamp 1554483974
transform 1 0 348 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_772
timestamp 1554483974
transform 1 0 348 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_1019
timestamp 1554483974
transform 1 0 380 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_743
timestamp 1554483974
transform 1 0 484 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_991
timestamp 1554483974
transform 1 0 484 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1020
timestamp 1554483974
transform 1 0 460 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_744
timestamp 1554483974
transform 1 0 516 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_745
timestamp 1554483974
transform 1 0 588 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_992
timestamp 1554483974
transform 1 0 516 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1021
timestamp 1554483974
transform 1 0 540 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_774
timestamp 1554483974
transform 1 0 588 0 1 295
box -3 -3 3 3
use M2_M1  M2_M1_985
timestamp 1554483974
transform 1 0 604 0 1 345
box -2 -2 2 2
use M3_M2  M3_M2_752
timestamp 1554483974
transform 1 0 604 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_993
timestamp 1554483974
transform 1 0 620 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_734
timestamp 1554483974
transform 1 0 636 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1022
timestamp 1554483974
transform 1 0 636 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1023
timestamp 1554483974
transform 1 0 660 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_986
timestamp 1554483974
transform 1 0 716 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_994
timestamp 1554483974
transform 1 0 700 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_753
timestamp 1554483974
transform 1 0 716 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_995
timestamp 1554483974
transform 1 0 724 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1024
timestamp 1554483974
transform 1 0 692 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_763
timestamp 1554483974
transform 1 0 700 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_764
timestamp 1554483974
transform 1 0 724 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1046
timestamp 1554483974
transform 1 0 724 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_754
timestamp 1554483974
transform 1 0 820 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1025
timestamp 1554483974
transform 1 0 820 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1047
timestamp 1554483974
transform 1 0 820 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1058
timestamp 1554483974
transform 1 0 812 0 1 305
box -2 -2 2 2
use M3_M2  M3_M2_775
timestamp 1554483974
transform 1 0 812 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_737
timestamp 1554483974
transform 1 0 916 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_738
timestamp 1554483974
transform 1 0 948 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_746
timestamp 1554483974
transform 1 0 924 0 1 345
box -3 -3 3 3
use M3_M2  M3_M2_747
timestamp 1554483974
transform 1 0 948 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_996
timestamp 1554483974
transform 1 0 916 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_755
timestamp 1554483974
transform 1 0 924 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_997
timestamp 1554483974
transform 1 0 932 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_998
timestamp 1554483974
transform 1 0 948 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1026
timestamp 1554483974
transform 1 0 924 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1027
timestamp 1554483974
transform 1 0 940 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_735
timestamp 1554483974
transform 1 0 964 0 1 365
box -3 -3 3 3
use M3_M2  M3_M2_776
timestamp 1554483974
transform 1 0 972 0 1 295
box -3 -3 3 3
use M3_M2  M3_M2_736
timestamp 1554483974
transform 1 0 1028 0 1 365
box -3 -3 3 3
use M2_M1  M2_M1_1028
timestamp 1554483974
transform 1 0 1028 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1048
timestamp 1554483974
transform 1 0 1020 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1059
timestamp 1554483974
transform 1 0 1036 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1060
timestamp 1554483974
transform 1 0 1052 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_1029
timestamp 1554483974
transform 1 0 1084 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1049
timestamp 1554483974
transform 1 0 1068 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1050
timestamp 1554483974
transform 1 0 1076 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1061
timestamp 1554483974
transform 1 0 1092 0 1 305
box -2 -2 2 2
use M2_M1  M2_M1_999
timestamp 1554483974
transform 1 0 1148 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1051
timestamp 1554483974
transform 1 0 1132 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_767
timestamp 1554483974
transform 1 0 1140 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1000
timestamp 1554483974
transform 1 0 1188 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_765
timestamp 1554483974
transform 1 0 1180 0 1 325
box -3 -3 3 3
use M2_M1  M2_M1_1001
timestamp 1554483974
transform 1 0 1212 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1030
timestamp 1554483974
transform 1 0 1204 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1052
timestamp 1554483974
transform 1 0 1180 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_766
timestamp 1554483974
transform 1 0 1212 0 1 325
box -3 -3 3 3
use M3_M2  M3_M2_768
timestamp 1554483974
transform 1 0 1204 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_748
timestamp 1554483974
transform 1 0 1244 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1002
timestamp 1554483974
transform 1 0 1244 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1003
timestamp 1554483974
transform 1 0 1252 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_749
timestamp 1554483974
transform 1 0 1292 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1004
timestamp 1554483974
transform 1 0 1276 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_756
timestamp 1554483974
transform 1 0 1284 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1005
timestamp 1554483974
transform 1 0 1300 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1031
timestamp 1554483974
transform 1 0 1284 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1032
timestamp 1554483974
transform 1 0 1292 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_769
timestamp 1554483974
transform 1 0 1284 0 1 315
box -3 -3 3 3
use M2_M1  M2_M1_1053
timestamp 1554483974
transform 1 0 1292 0 1 315
box -2 -2 2 2
use M3_M2  M3_M2_770
timestamp 1554483974
transform 1 0 1300 0 1 315
box -3 -3 3 3
use M3_M2  M3_M2_773
timestamp 1554483974
transform 1 0 1292 0 1 305
box -3 -3 3 3
use M2_M1  M2_M1_987
timestamp 1554483974
transform 1 0 1372 0 1 345
box -2 -2 2 2
use M2_M1  M2_M1_1006
timestamp 1554483974
transform 1 0 1364 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_757
timestamp 1554483974
transform 1 0 1372 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1033
timestamp 1554483974
transform 1 0 1396 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_739
timestamp 1554483974
transform 1 0 1436 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_740
timestamp 1554483974
transform 1 0 1452 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1007
timestamp 1554483974
transform 1 0 1436 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1034
timestamp 1554483974
transform 1 0 1444 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1054
timestamp 1554483974
transform 1 0 1444 0 1 315
box -2 -2 2 2
use M2_M1  M2_M1_1008
timestamp 1554483974
transform 1 0 1476 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_741
timestamp 1554483974
transform 1 0 1492 0 1 355
box -3 -3 3 3
use M2_M1  M2_M1_1009
timestamp 1554483974
transform 1 0 1492 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_758
timestamp 1554483974
transform 1 0 1508 0 1 335
box -3 -3 3 3
use M3_M2  M3_M2_759
timestamp 1554483974
transform 1 0 1524 0 1 335
box -3 -3 3 3
use M2_M1  M2_M1_1035
timestamp 1554483974
transform 1 0 1500 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1036
timestamp 1554483974
transform 1 0 1524 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1010
timestamp 1554483974
transform 1 0 1540 0 1 335
box -2 -2 2 2
use M3_M2  M3_M2_742
timestamp 1554483974
transform 1 0 1588 0 1 355
box -3 -3 3 3
use M3_M2  M3_M2_750
timestamp 1554483974
transform 1 0 1572 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1011
timestamp 1554483974
transform 1 0 1580 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1012
timestamp 1554483974
transform 1 0 1596 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1037
timestamp 1554483974
transform 1 0 1572 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1038
timestamp 1554483974
transform 1 0 1588 0 1 325
box -2 -2 2 2
use M3_M2  M3_M2_751
timestamp 1554483974
transform 1 0 1676 0 1 345
box -3 -3 3 3
use M2_M1  M2_M1_1013
timestamp 1554483974
transform 1 0 1660 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1014
timestamp 1554483974
transform 1 0 1676 0 1 335
box -2 -2 2 2
use M2_M1  M2_M1_1039
timestamp 1554483974
transform 1 0 1652 0 1 325
box -2 -2 2 2
use M2_M1  M2_M1_1040
timestamp 1554483974
transform 1 0 1668 0 1 325
box -2 -2 2 2
use UART_VIA1  UART_VIA1_26
timestamp 1554483974
transform 1 0 24 0 1 270
box -10 -3 10 3
use FILL  FILL_858
timestamp 1554483974
transform 1 0 72 0 -1 370
box -8 -3 16 105
use FILL  FILL_860
timestamp 1554483974
transform 1 0 80 0 -1 370
box -8 -3 16 105
use FILL  FILL_862
timestamp 1554483974
transform 1 0 88 0 -1 370
box -8 -3 16 105
use FILL  FILL_865
timestamp 1554483974
transform 1 0 96 0 -1 370
box -8 -3 16 105
use FILL  FILL_866
timestamp 1554483974
transform 1 0 104 0 -1 370
box -8 -3 16 105
use FILL  FILL_867
timestamp 1554483974
transform 1 0 112 0 -1 370
box -8 -3 16 105
use FILL  FILL_868
timestamp 1554483974
transform 1 0 120 0 -1 370
box -8 -3 16 105
use FILL  FILL_869
timestamp 1554483974
transform 1 0 128 0 -1 370
box -8 -3 16 105
use FILL  FILL_870
timestamp 1554483974
transform 1 0 136 0 -1 370
box -8 -3 16 105
use FILL  FILL_872
timestamp 1554483974
transform 1 0 144 0 -1 370
box -8 -3 16 105
use FILL  FILL_874
timestamp 1554483974
transform 1 0 152 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_12
timestamp 1554483974
transform 1 0 160 0 -1 370
box -8 -3 40 105
use FILL  FILL_878
timestamp 1554483974
transform 1 0 192 0 -1 370
box -8 -3 16 105
use FILL  FILL_879
timestamp 1554483974
transform 1 0 200 0 -1 370
box -8 -3 16 105
use FILL  FILL_880
timestamp 1554483974
transform 1 0 208 0 -1 370
box -8 -3 16 105
use FILL  FILL_882
timestamp 1554483974
transform 1 0 216 0 -1 370
box -8 -3 16 105
use FILL  FILL_884
timestamp 1554483974
transform 1 0 224 0 -1 370
box -8 -3 16 105
use FILL  FILL_889
timestamp 1554483974
transform 1 0 232 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_13
timestamp 1554483974
transform -1 0 272 0 -1 370
box -8 -3 40 105
use FILL  FILL_890
timestamp 1554483974
transform 1 0 272 0 -1 370
box -8 -3 16 105
use FILL  FILL_892
timestamp 1554483974
transform 1 0 280 0 -1 370
box -8 -3 16 105
use FILL  FILL_894
timestamp 1554483974
transform 1 0 288 0 -1 370
box -8 -3 16 105
use FILL  FILL_896
timestamp 1554483974
transform 1 0 296 0 -1 370
box -8 -3 16 105
use FILL  FILL_898
timestamp 1554483974
transform 1 0 304 0 -1 370
box -8 -3 16 105
use FILL  FILL_900
timestamp 1554483974
transform 1 0 312 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_18
timestamp 1554483974
transform 1 0 320 0 -1 370
box -8 -3 46 105
use FILL  FILL_902
timestamp 1554483974
transform 1 0 360 0 -1 370
box -8 -3 16 105
use FILL  FILL_904
timestamp 1554483974
transform 1 0 368 0 -1 370
box -8 -3 16 105
use FILL  FILL_906
timestamp 1554483974
transform 1 0 376 0 -1 370
box -8 -3 16 105
use FILL  FILL_908
timestamp 1554483974
transform 1 0 384 0 -1 370
box -8 -3 16 105
use FILL  FILL_913
timestamp 1554483974
transform 1 0 392 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_46
timestamp 1554483974
transform -1 0 496 0 -1 370
box -8 -3 104 105
use FILL  FILL_914
timestamp 1554483974
transform 1 0 496 0 -1 370
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_47
timestamp 1554483974
transform 1 0 504 0 -1 370
box -8 -3 104 105
use FILL  FILL_915
timestamp 1554483974
transform 1 0 600 0 -1 370
box -8 -3 16 105
use FILL  FILL_916
timestamp 1554483974
transform 1 0 608 0 -1 370
box -8 -3 16 105
use FILL  FILL_917
timestamp 1554483974
transform 1 0 616 0 -1 370
box -8 -3 16 105
use FILL  FILL_918
timestamp 1554483974
transform 1 0 624 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_13
timestamp 1554483974
transform 1 0 632 0 -1 370
box -8 -3 32 105
use FILL  FILL_919
timestamp 1554483974
transform 1 0 656 0 -1 370
box -8 -3 16 105
use FILL  FILL_920
timestamp 1554483974
transform 1 0 664 0 -1 370
box -8 -3 16 105
use FILL  FILL_921
timestamp 1554483974
transform 1 0 672 0 -1 370
box -8 -3 16 105
use FILL  FILL_923
timestamp 1554483974
transform 1 0 680 0 -1 370
box -8 -3 16 105
use AOI21X1  AOI21X1_3
timestamp 1554483974
transform 1 0 688 0 -1 370
box -7 -3 39 105
use FILL  FILL_927
timestamp 1554483974
transform 1 0 720 0 -1 370
box -8 -3 16 105
use FILL  FILL_928
timestamp 1554483974
transform 1 0 728 0 -1 370
box -8 -3 16 105
use FILL  FILL_929
timestamp 1554483974
transform 1 0 736 0 -1 370
box -8 -3 16 105
use FILL  FILL_930
timestamp 1554483974
transform 1 0 744 0 -1 370
box -8 -3 16 105
use FILL  FILL_931
timestamp 1554483974
transform 1 0 752 0 -1 370
box -8 -3 16 105
use FILL  FILL_932
timestamp 1554483974
transform 1 0 760 0 -1 370
box -8 -3 16 105
use FILL  FILL_933
timestamp 1554483974
transform 1 0 768 0 -1 370
box -8 -3 16 105
use FILL  FILL_934
timestamp 1554483974
transform 1 0 776 0 -1 370
box -8 -3 16 105
use FILL  FILL_935
timestamp 1554483974
transform 1 0 784 0 -1 370
box -8 -3 16 105
use FILL  FILL_936
timestamp 1554483974
transform 1 0 792 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_14
timestamp 1554483974
transform -1 0 832 0 -1 370
box -8 -3 40 105
use FILL  FILL_937
timestamp 1554483974
transform 1 0 832 0 -1 370
box -8 -3 16 105
use FILL  FILL_938
timestamp 1554483974
transform 1 0 840 0 -1 370
box -8 -3 16 105
use FILL  FILL_939
timestamp 1554483974
transform 1 0 848 0 -1 370
box -8 -3 16 105
use FILL  FILL_940
timestamp 1554483974
transform 1 0 856 0 -1 370
box -8 -3 16 105
use FILL  FILL_941
timestamp 1554483974
transform 1 0 864 0 -1 370
box -8 -3 16 105
use FILL  FILL_943
timestamp 1554483974
transform 1 0 872 0 -1 370
box -8 -3 16 105
use FILL  FILL_945
timestamp 1554483974
transform 1 0 880 0 -1 370
box -8 -3 16 105
use FILL  FILL_947
timestamp 1554483974
transform 1 0 888 0 -1 370
box -8 -3 16 105
use FILL  FILL_949
timestamp 1554483974
transform 1 0 896 0 -1 370
box -8 -3 16 105
use FILL  FILL_953
timestamp 1554483974
transform 1 0 904 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_19
timestamp 1554483974
transform -1 0 952 0 -1 370
box -8 -3 46 105
use FILL  FILL_954
timestamp 1554483974
transform 1 0 952 0 -1 370
box -8 -3 16 105
use FILL  FILL_956
timestamp 1554483974
transform 1 0 960 0 -1 370
box -8 -3 16 105
use FILL  FILL_957
timestamp 1554483974
transform 1 0 968 0 -1 370
box -8 -3 16 105
use FILL  FILL_958
timestamp 1554483974
transform 1 0 976 0 -1 370
box -8 -3 16 105
use FILL  FILL_960
timestamp 1554483974
transform 1 0 984 0 -1 370
box -8 -3 16 105
use FILL  FILL_962
timestamp 1554483974
transform 1 0 992 0 -1 370
box -8 -3 16 105
use FILL  FILL_966
timestamp 1554483974
transform 1 0 1000 0 -1 370
box -8 -3 16 105
use FILL  FILL_967
timestamp 1554483974
transform 1 0 1008 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_16
timestamp 1554483974
transform 1 0 1016 0 -1 370
box -8 -3 40 105
use FILL  FILL_968
timestamp 1554483974
transform 1 0 1048 0 -1 370
box -8 -3 16 105
use FILL  FILL_970
timestamp 1554483974
transform 1 0 1056 0 -1 370
box -8 -3 16 105
use FILL  FILL_972
timestamp 1554483974
transform 1 0 1064 0 -1 370
box -8 -3 16 105
use NAND3X1  NAND3X1_17
timestamp 1554483974
transform 1 0 1072 0 -1 370
box -8 -3 40 105
use FILL  FILL_976
timestamp 1554483974
transform 1 0 1104 0 -1 370
box -8 -3 16 105
use FILL  FILL_989
timestamp 1554483974
transform 1 0 1112 0 -1 370
box -8 -3 16 105
use FILL  FILL_990
timestamp 1554483974
transform 1 0 1120 0 -1 370
box -8 -3 16 105
use FILL  FILL_991
timestamp 1554483974
transform 1 0 1128 0 -1 370
box -8 -3 16 105
use FILL  FILL_992
timestamp 1554483974
transform 1 0 1136 0 -1 370
box -8 -3 16 105
use FILL  FILL_993
timestamp 1554483974
transform 1 0 1144 0 -1 370
box -8 -3 16 105
use FILL  FILL_994
timestamp 1554483974
transform 1 0 1152 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_51
timestamp 1554483974
transform 1 0 1160 0 -1 370
box -8 -3 32 105
use OAI21X1  OAI21X1_38
timestamp 1554483974
transform -1 0 1216 0 -1 370
box -8 -3 34 105
use FILL  FILL_995
timestamp 1554483974
transform 1 0 1216 0 -1 370
box -8 -3 16 105
use FILL  FILL_996
timestamp 1554483974
transform 1 0 1224 0 -1 370
box -8 -3 16 105
use FILL  FILL_997
timestamp 1554483974
transform 1 0 1232 0 -1 370
box -8 -3 16 105
use FILL  FILL_998
timestamp 1554483974
transform 1 0 1240 0 -1 370
box -8 -3 16 105
use FILL  FILL_999
timestamp 1554483974
transform 1 0 1248 0 -1 370
box -8 -3 16 105
use FILL  FILL_1000
timestamp 1554483974
transform 1 0 1256 0 -1 370
box -8 -3 16 105
use FILL  FILL_1001
timestamp 1554483974
transform 1 0 1264 0 -1 370
box -8 -3 16 105
use NAND2X1  NAND2X1_52
timestamp 1554483974
transform 1 0 1272 0 -1 370
box -8 -3 32 105
use INVX2  INVX2_69
timestamp 1554483974
transform 1 0 1296 0 -1 370
box -9 -3 26 105
use FILL  FILL_1002
timestamp 1554483974
transform 1 0 1312 0 -1 370
box -8 -3 16 105
use FILL  FILL_1004
timestamp 1554483974
transform 1 0 1320 0 -1 370
box -8 -3 16 105
use FILL  FILL_1008
timestamp 1554483974
transform 1 0 1328 0 -1 370
box -8 -3 16 105
use FILL  FILL_1009
timestamp 1554483974
transform 1 0 1336 0 -1 370
box -8 -3 16 105
use FILL  FILL_1010
timestamp 1554483974
transform 1 0 1344 0 -1 370
box -8 -3 16 105
use NOR2X1  NOR2X1_14
timestamp 1554483974
transform -1 0 1376 0 -1 370
box -8 -3 32 105
use FILL  FILL_1011
timestamp 1554483974
transform 1 0 1376 0 -1 370
box -8 -3 16 105
use FILL  FILL_1013
timestamp 1554483974
transform 1 0 1384 0 -1 370
box -8 -3 16 105
use FILL  FILL_1015
timestamp 1554483974
transform 1 0 1392 0 -1 370
box -8 -3 16 105
use FILL  FILL_1017
timestamp 1554483974
transform 1 0 1400 0 -1 370
box -8 -3 16 105
use FILL  FILL_1019
timestamp 1554483974
transform 1 0 1408 0 -1 370
box -8 -3 16 105
use FILL  FILL_1023
timestamp 1554483974
transform 1 0 1416 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_70
timestamp 1554483974
transform -1 0 1440 0 -1 370
box -9 -3 26 105
use NAND2X1  NAND2X1_53
timestamp 1554483974
transform -1 0 1464 0 -1 370
box -8 -3 32 105
use FILL  FILL_1024
timestamp 1554483974
transform 1 0 1464 0 -1 370
box -8 -3 16 105
use FILL  FILL_1026
timestamp 1554483974
transform 1 0 1472 0 -1 370
box -8 -3 16 105
use FILL  FILL_1028
timestamp 1554483974
transform 1 0 1480 0 -1 370
box -8 -3 16 105
use FILL  FILL_1030
timestamp 1554483974
transform 1 0 1488 0 -1 370
box -8 -3 16 105
use AOI21X1  AOI21X1_4
timestamp 1554483974
transform 1 0 1496 0 -1 370
box -7 -3 39 105
use FILL  FILL_1031
timestamp 1554483974
transform 1 0 1528 0 -1 370
box -8 -3 16 105
use FILL  FILL_1033
timestamp 1554483974
transform 1 0 1536 0 -1 370
box -8 -3 16 105
use FILL  FILL_1035
timestamp 1554483974
transform 1 0 1544 0 -1 370
box -8 -3 16 105
use FILL  FILL_1037
timestamp 1554483974
transform 1 0 1552 0 -1 370
box -8 -3 16 105
use INVX2  INVX2_73
timestamp 1554483974
transform 1 0 1560 0 -1 370
box -9 -3 26 105
use NAND2X1  NAND2X1_55
timestamp 1554483974
transform 1 0 1576 0 -1 370
box -8 -3 32 105
use FILL  FILL_1046
timestamp 1554483974
transform 1 0 1600 0 -1 370
box -8 -3 16 105
use FILL  FILL_1047
timestamp 1554483974
transform 1 0 1608 0 -1 370
box -8 -3 16 105
use FILL  FILL_1048
timestamp 1554483974
transform 1 0 1616 0 -1 370
box -8 -3 16 105
use FILL  FILL_1049
timestamp 1554483974
transform 1 0 1624 0 -1 370
box -8 -3 16 105
use FILL  FILL_1050
timestamp 1554483974
transform 1 0 1632 0 -1 370
box -8 -3 16 105
use OAI22X1  OAI22X1_22
timestamp 1554483974
transform -1 0 1680 0 -1 370
box -8 -3 46 105
use FILL  FILL_1051
timestamp 1554483974
transform 1 0 1680 0 -1 370
box -8 -3 16 105
use FILL  FILL_1052
timestamp 1554483974
transform 1 0 1688 0 -1 370
box -8 -3 16 105
use FILL  FILL_1053
timestamp 1554483974
transform 1 0 1696 0 -1 370
box -8 -3 16 105
use FILL  FILL_1054
timestamp 1554483974
transform 1 0 1704 0 -1 370
box -8 -3 16 105
use FILL  FILL_1055
timestamp 1554483974
transform 1 0 1712 0 -1 370
box -8 -3 16 105
use FILL  FILL_1056
timestamp 1554483974
transform 1 0 1720 0 -1 370
box -8 -3 16 105
use FILL  FILL_1057
timestamp 1554483974
transform 1 0 1728 0 -1 370
box -8 -3 16 105
use FILL  FILL_1058
timestamp 1554483974
transform 1 0 1736 0 -1 370
box -8 -3 16 105
use FILL  FILL_1059
timestamp 1554483974
transform 1 0 1744 0 -1 370
box -8 -3 16 105
use FILL  FILL_1060
timestamp 1554483974
transform 1 0 1752 0 -1 370
box -8 -3 16 105
use FILL  FILL_1061
timestamp 1554483974
transform 1 0 1760 0 -1 370
box -8 -3 16 105
use FILL  FILL_1062
timestamp 1554483974
transform 1 0 1768 0 -1 370
box -8 -3 16 105
use UART_VIA1  UART_VIA1_27
timestamp 1554483974
transform 1 0 1825 0 1 270
box -10 -3 10 3
use M2_M1  M2_M1_1109
timestamp 1554483974
transform 1 0 76 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1067
timestamp 1554483974
transform 1 0 108 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_800
timestamp 1554483974
transform 1 0 132 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1110
timestamp 1554483974
transform 1 0 132 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1080
timestamp 1554483974
transform 1 0 164 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1081
timestamp 1554483974
transform 1 0 172 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1111
timestamp 1554483974
transform 1 0 220 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_820
timestamp 1554483974
transform 1 0 220 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_801
timestamp 1554483974
transform 1 0 236 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1112
timestamp 1554483974
transform 1 0 236 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_782
timestamp 1554483974
transform 1 0 260 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_783
timestamp 1554483974
transform 1 0 364 0 1 235
box -3 -3 3 3
use M3_M2  M3_M2_790
timestamp 1554483974
transform 1 0 348 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1068
timestamp 1554483974
transform 1 0 364 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1082
timestamp 1554483974
transform 1 0 260 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1083
timestamp 1554483974
transform 1 0 268 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1084
timestamp 1554483974
transform 1 0 324 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1113
timestamp 1554483974
transform 1 0 348 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_821
timestamp 1554483974
transform 1 0 268 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1114
timestamp 1554483974
transform 1 0 380 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1135
timestamp 1554483974
transform 1 0 396 0 1 195
box -2 -2 2 2
use M2_M1  M2_M1_1085
timestamp 1554483974
transform 1 0 436 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1086
timestamp 1554483974
transform 1 0 452 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1115
timestamp 1554483974
transform 1 0 460 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1087
timestamp 1554483974
transform 1 0 532 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_812
timestamp 1554483974
transform 1 0 532 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1136
timestamp 1554483974
transform 1 0 532 0 1 195
box -2 -2 2 2
use M3_M2  M3_M2_791
timestamp 1554483974
transform 1 0 556 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1088
timestamp 1554483974
transform 1 0 556 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_813
timestamp 1554483974
transform 1 0 604 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_802
timestamp 1554483974
transform 1 0 628 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1116
timestamp 1554483974
transform 1 0 628 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1117
timestamp 1554483974
transform 1 0 636 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_822
timestamp 1554483974
transform 1 0 636 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1089
timestamp 1554483974
transform 1 0 660 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_823
timestamp 1554483974
transform 1 0 660 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_784
timestamp 1554483974
transform 1 0 684 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1062
timestamp 1554483974
transform 1 0 700 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_785
timestamp 1554483974
transform 1 0 708 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1069
timestamp 1554483974
transform 1 0 684 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1070
timestamp 1554483974
transform 1 0 692 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1090
timestamp 1554483974
transform 1 0 708 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1071
timestamp 1554483974
transform 1 0 740 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1063
timestamp 1554483974
transform 1 0 820 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_792
timestamp 1554483974
transform 1 0 812 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1072
timestamp 1554483974
transform 1 0 828 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1091
timestamp 1554483974
transform 1 0 812 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_803
timestamp 1554483974
transform 1 0 828 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_814
timestamp 1554483974
transform 1 0 820 0 1 205
box -3 -3 3 3
use M3_M2  M3_M2_793
timestamp 1554483974
transform 1 0 924 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_786
timestamp 1554483974
transform 1 0 956 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1092
timestamp 1554483974
transform 1 0 924 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_804
timestamp 1554483974
transform 1 0 948 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1093
timestamp 1554483974
transform 1 0 956 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1118
timestamp 1554483974
transform 1 0 916 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1119
timestamp 1554483974
transform 1 0 932 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1120
timestamp 1554483974
transform 1 0 948 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1121
timestamp 1554483974
transform 1 0 956 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_824
timestamp 1554483974
transform 1 0 916 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_825
timestamp 1554483974
transform 1 0 956 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_777
timestamp 1554483974
transform 1 0 1020 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_779
timestamp 1554483974
transform 1 0 1020 0 1 245
box -3 -3 3 3
use M3_M2  M3_M2_794
timestamp 1554483974
transform 1 0 1036 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_778
timestamp 1554483974
transform 1 0 1060 0 1 255
box -3 -3 3 3
use M3_M2  M3_M2_787
timestamp 1554483974
transform 1 0 1052 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1064
timestamp 1554483974
transform 1 0 1060 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1073
timestamp 1554483974
transform 1 0 1052 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1094
timestamp 1554483974
transform 1 0 1020 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1095
timestamp 1554483974
transform 1 0 1036 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_805
timestamp 1554483974
transform 1 0 1044 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1122
timestamp 1554483974
transform 1 0 1028 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1123
timestamp 1554483974
transform 1 0 1044 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_795
timestamp 1554483974
transform 1 0 1084 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1096
timestamp 1554483974
transform 1 0 1084 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_780
timestamp 1554483974
transform 1 0 1132 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_1074
timestamp 1554483974
transform 1 0 1132 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_815
timestamp 1554483974
transform 1 0 1124 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1097
timestamp 1554483974
transform 1 0 1148 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1098
timestamp 1554483974
transform 1 0 1188 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_816
timestamp 1554483974
transform 1 0 1204 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1124
timestamp 1554483974
transform 1 0 1228 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_781
timestamp 1554483974
transform 1 0 1252 0 1 245
box -3 -3 3 3
use M2_M1  M2_M1_1099
timestamp 1554483974
transform 1 0 1244 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_817
timestamp 1554483974
transform 1 0 1244 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1125
timestamp 1554483974
transform 1 0 1284 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_826
timestamp 1554483974
transform 1 0 1284 0 1 195
box -3 -3 3 3
use M2_M1  M2_M1_1126
timestamp 1554483974
transform 1 0 1308 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_788
timestamp 1554483974
transform 1 0 1364 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1075
timestamp 1554483974
transform 1 0 1364 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1065
timestamp 1554483974
transform 1 0 1380 0 1 235
box -2 -2 2 2
use M2_M1  M2_M1_1100
timestamp 1554483974
transform 1 0 1364 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_806
timestamp 1554483974
transform 1 0 1372 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1076
timestamp 1554483974
transform 1 0 1396 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1066
timestamp 1554483974
transform 1 0 1460 0 1 235
box -2 -2 2 2
use M3_M2  M3_M2_796
timestamp 1554483974
transform 1 0 1460 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1101
timestamp 1554483974
transform 1 0 1452 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_807
timestamp 1554483974
transform 1 0 1468 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1077
timestamp 1554483974
transform 1 0 1492 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_808
timestamp 1554483974
transform 1 0 1484 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_818
timestamp 1554483974
transform 1 0 1476 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1127
timestamp 1554483974
transform 1 0 1484 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1102
timestamp 1554483974
transform 1 0 1508 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_797
timestamp 1554483974
transform 1 0 1532 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1103
timestamp 1554483974
transform 1 0 1532 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1078
timestamp 1554483974
transform 1 0 1548 0 1 225
box -2 -2 2 2
use M2_M1  M2_M1_1128
timestamp 1554483974
transform 1 0 1540 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_827
timestamp 1554483974
transform 1 0 1548 0 1 195
box -3 -3 3 3
use M3_M2  M3_M2_789
timestamp 1554483974
transform 1 0 1588 0 1 235
box -3 -3 3 3
use M2_M1  M2_M1_1129
timestamp 1554483974
transform 1 0 1588 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1130
timestamp 1554483974
transform 1 0 1620 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1079
timestamp 1554483974
transform 1 0 1636 0 1 225
box -2 -2 2 2
use M3_M2  M3_M2_798
timestamp 1554483974
transform 1 0 1660 0 1 225
box -3 -3 3 3
use M3_M2  M3_M2_809
timestamp 1554483974
transform 1 0 1636 0 1 215
box -3 -3 3 3
use M3_M2  M3_M2_799
timestamp 1554483974
transform 1 0 1716 0 1 225
box -3 -3 3 3
use M2_M1  M2_M1_1104
timestamp 1554483974
transform 1 0 1644 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1105
timestamp 1554483974
transform 1 0 1652 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1106
timestamp 1554483974
transform 1 0 1668 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_810
timestamp 1554483974
transform 1 0 1676 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1107
timestamp 1554483974
transform 1 0 1716 0 1 215
box -2 -2 2 2
use M3_M2  M3_M2_811
timestamp 1554483974
transform 1 0 1772 0 1 215
box -3 -3 3 3
use M2_M1  M2_M1_1108
timestamp 1554483974
transform 1 0 1780 0 1 215
box -2 -2 2 2
use M2_M1  M2_M1_1131
timestamp 1554483974
transform 1 0 1644 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_819
timestamp 1554483974
transform 1 0 1652 0 1 205
box -3 -3 3 3
use M2_M1  M2_M1_1132
timestamp 1554483974
transform 1 0 1660 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1133
timestamp 1554483974
transform 1 0 1676 0 1 205
box -2 -2 2 2
use M2_M1  M2_M1_1134
timestamp 1554483974
transform 1 0 1692 0 1 205
box -2 -2 2 2
use M3_M2  M3_M2_828
timestamp 1554483974
transform 1 0 1644 0 1 195
box -3 -3 3 3
use UART_VIA1  UART_VIA1_28
timestamp 1554483974
transform 1 0 48 0 1 170
box -10 -3 10 3
use FILL  FILL_1063
timestamp 1554483974
transform 1 0 72 0 1 170
box -8 -3 16 105
use FILL  FILL_1065
timestamp 1554483974
transform 1 0 80 0 1 170
box -8 -3 16 105
use FILL  FILL_1067
timestamp 1554483974
transform 1 0 88 0 1 170
box -8 -3 16 105
use FILL  FILL_1069
timestamp 1554483974
transform 1 0 96 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_40
timestamp 1554483974
transform -1 0 136 0 1 170
box -8 -3 34 105
use FILL  FILL_1070
timestamp 1554483974
transform 1 0 136 0 1 170
box -8 -3 16 105
use FILL  FILL_1077
timestamp 1554483974
transform 1 0 144 0 1 170
box -8 -3 16 105
use FILL  FILL_1079
timestamp 1554483974
transform 1 0 152 0 1 170
box -8 -3 16 105
use FILL  FILL_1080
timestamp 1554483974
transform 1 0 160 0 1 170
box -8 -3 16 105
use FILL  FILL_1081
timestamp 1554483974
transform 1 0 168 0 1 170
box -8 -3 16 105
use FILL  FILL_1082
timestamp 1554483974
transform 1 0 176 0 1 170
box -8 -3 16 105
use FILL  FILL_1085
timestamp 1554483974
transform 1 0 184 0 1 170
box -8 -3 16 105
use FILL  FILL_1087
timestamp 1554483974
transform 1 0 192 0 1 170
box -8 -3 16 105
use FILL  FILL_1089
timestamp 1554483974
transform 1 0 200 0 1 170
box -8 -3 16 105
use INVX2  INVX2_75
timestamp 1554483974
transform -1 0 224 0 1 170
box -9 -3 26 105
use FILL  FILL_1090
timestamp 1554483974
transform 1 0 224 0 1 170
box -8 -3 16 105
use FILL  FILL_1091
timestamp 1554483974
transform 1 0 232 0 1 170
box -8 -3 16 105
use FILL  FILL_1092
timestamp 1554483974
transform 1 0 240 0 1 170
box -8 -3 16 105
use INVX2  INVX2_76
timestamp 1554483974
transform 1 0 248 0 1 170
box -9 -3 26 105
use DFFNEGX1  DFFNEGX1_50
timestamp 1554483974
transform -1 0 360 0 1 170
box -8 -3 104 105
use NAND2X1  NAND2X1_56
timestamp 1554483974
transform -1 0 384 0 1 170
box -8 -3 32 105
use FILL  FILL_1095
timestamp 1554483974
transform 1 0 384 0 1 170
box -8 -3 16 105
use FILL  FILL_1110
timestamp 1554483974
transform 1 0 392 0 1 170
box -8 -3 16 105
use FILL  FILL_1112
timestamp 1554483974
transform 1 0 400 0 1 170
box -8 -3 16 105
use FILL  FILL_1114
timestamp 1554483974
transform 1 0 408 0 1 170
box -8 -3 16 105
use FILL  FILL_1116
timestamp 1554483974
transform 1 0 416 0 1 170
box -8 -3 16 105
use FILL  FILL_1118
timestamp 1554483974
transform 1 0 424 0 1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_15
timestamp 1554483974
transform 1 0 432 0 1 170
box -8 -3 32 105
use FILL  FILL_1120
timestamp 1554483974
transform 1 0 456 0 1 170
box -8 -3 16 105
use FILL  FILL_1125
timestamp 1554483974
transform 1 0 464 0 1 170
box -8 -3 16 105
use FILL  FILL_1127
timestamp 1554483974
transform 1 0 472 0 1 170
box -8 -3 16 105
use FILL  FILL_1129
timestamp 1554483974
transform 1 0 480 0 1 170
box -8 -3 16 105
use FILL  FILL_1130
timestamp 1554483974
transform 1 0 488 0 1 170
box -8 -3 16 105
use FILL  FILL_1131
timestamp 1554483974
transform 1 0 496 0 1 170
box -8 -3 16 105
use FILL  FILL_1133
timestamp 1554483974
transform 1 0 504 0 1 170
box -8 -3 16 105
use FILL  FILL_1135
timestamp 1554483974
transform 1 0 512 0 1 170
box -8 -3 16 105
use FILL  FILL_1137
timestamp 1554483974
transform 1 0 520 0 1 170
box -8 -3 16 105
use AOI21X1  AOI21X1_5
timestamp 1554483974
transform -1 0 560 0 1 170
box -7 -3 39 105
use FILL  FILL_1138
timestamp 1554483974
transform 1 0 560 0 1 170
box -8 -3 16 105
use FILL  FILL_1139
timestamp 1554483974
transform 1 0 568 0 1 170
box -8 -3 16 105
use FILL  FILL_1140
timestamp 1554483974
transform 1 0 576 0 1 170
box -8 -3 16 105
use FILL  FILL_1141
timestamp 1554483974
transform 1 0 584 0 1 170
box -8 -3 16 105
use FILL  FILL_1147
timestamp 1554483974
transform 1 0 592 0 1 170
box -8 -3 16 105
use FILL  FILL_1149
timestamp 1554483974
transform 1 0 600 0 1 170
box -8 -3 16 105
use FILL  FILL_1151
timestamp 1554483974
transform 1 0 608 0 1 170
box -8 -3 16 105
use FILL  FILL_1153
timestamp 1554483974
transform 1 0 616 0 1 170
box -8 -3 16 105
use FILL  FILL_1154
timestamp 1554483974
transform 1 0 624 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_57
timestamp 1554483974
transform 1 0 632 0 1 170
box -8 -3 32 105
use FILL  FILL_1155
timestamp 1554483974
transform 1 0 656 0 1 170
box -8 -3 16 105
use FILL  FILL_1156
timestamp 1554483974
transform 1 0 664 0 1 170
box -8 -3 16 105
use FILL  FILL_1157
timestamp 1554483974
transform 1 0 672 0 1 170
box -8 -3 16 105
use FILL  FILL_1158
timestamp 1554483974
transform 1 0 680 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_20
timestamp 1554483974
transform -1 0 720 0 1 170
box -8 -3 40 105
use FILL  FILL_1159
timestamp 1554483974
transform 1 0 720 0 1 170
box -8 -3 16 105
use FILL  FILL_1166
timestamp 1554483974
transform 1 0 728 0 1 170
box -8 -3 16 105
use FILL  FILL_1168
timestamp 1554483974
transform 1 0 736 0 1 170
box -8 -3 16 105
use FILL  FILL_1170
timestamp 1554483974
transform 1 0 744 0 1 170
box -8 -3 16 105
use FILL  FILL_1171
timestamp 1554483974
transform 1 0 752 0 1 170
box -8 -3 16 105
use FILL  FILL_1172
timestamp 1554483974
transform 1 0 760 0 1 170
box -8 -3 16 105
use FILL  FILL_1174
timestamp 1554483974
transform 1 0 768 0 1 170
box -8 -3 16 105
use FILL  FILL_1176
timestamp 1554483974
transform 1 0 776 0 1 170
box -8 -3 16 105
use FILL  FILL_1178
timestamp 1554483974
transform 1 0 784 0 1 170
box -8 -3 16 105
use FILL  FILL_1180
timestamp 1554483974
transform 1 0 792 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_22
timestamp 1554483974
transform 1 0 800 0 1 170
box -8 -3 40 105
use FILL  FILL_1182
timestamp 1554483974
transform 1 0 832 0 1 170
box -8 -3 16 105
use FILL  FILL_1186
timestamp 1554483974
transform 1 0 840 0 1 170
box -8 -3 16 105
use FILL  FILL_1188
timestamp 1554483974
transform 1 0 848 0 1 170
box -8 -3 16 105
use FILL  FILL_1190
timestamp 1554483974
transform 1 0 856 0 1 170
box -8 -3 16 105
use FILL  FILL_1192
timestamp 1554483974
transform 1 0 864 0 1 170
box -8 -3 16 105
use FILL  FILL_1193
timestamp 1554483974
transform 1 0 872 0 1 170
box -8 -3 16 105
use FILL  FILL_1194
timestamp 1554483974
transform 1 0 880 0 1 170
box -8 -3 16 105
use FILL  FILL_1195
timestamp 1554483974
transform 1 0 888 0 1 170
box -8 -3 16 105
use FILL  FILL_1196
timestamp 1554483974
transform 1 0 896 0 1 170
box -8 -3 16 105
use FILL  FILL_1197
timestamp 1554483974
transform 1 0 904 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_23
timestamp 1554483974
transform -1 0 952 0 1 170
box -8 -3 46 105
use FILL  FILL_1198
timestamp 1554483974
transform 1 0 952 0 1 170
box -8 -3 16 105
use FILL  FILL_1199
timestamp 1554483974
transform 1 0 960 0 1 170
box -8 -3 16 105
use FILL  FILL_1200
timestamp 1554483974
transform 1 0 968 0 1 170
box -8 -3 16 105
use FILL  FILL_1203
timestamp 1554483974
transform 1 0 976 0 1 170
box -8 -3 16 105
use FILL  FILL_1204
timestamp 1554483974
transform 1 0 984 0 1 170
box -8 -3 16 105
use FILL  FILL_1205
timestamp 1554483974
transform 1 0 992 0 1 170
box -8 -3 16 105
use FILL  FILL_1207
timestamp 1554483974
transform 1 0 1000 0 1 170
box -8 -3 16 105
use OAI22X1  OAI22X1_24
timestamp 1554483974
transform -1 0 1048 0 1 170
box -8 -3 46 105
use FILL  FILL_1208
timestamp 1554483974
transform 1 0 1048 0 1 170
box -8 -3 16 105
use FILL  FILL_1209
timestamp 1554483974
transform 1 0 1056 0 1 170
box -8 -3 16 105
use FILL  FILL_1210
timestamp 1554483974
transform 1 0 1064 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_23
timestamp 1554483974
transform 1 0 1072 0 1 170
box -8 -3 40 105
use FILL  FILL_1211
timestamp 1554483974
transform 1 0 1104 0 1 170
box -8 -3 16 105
use FILL  FILL_1212
timestamp 1554483974
transform 1 0 1112 0 1 170
box -8 -3 16 105
use FILL  FILL_1213
timestamp 1554483974
transform 1 0 1120 0 1 170
box -8 -3 16 105
use FILL  FILL_1218
timestamp 1554483974
transform 1 0 1128 0 1 170
box -8 -3 16 105
use FILL  FILL_1220
timestamp 1554483974
transform 1 0 1136 0 1 170
box -8 -3 16 105
use DFFNEGX1  DFFNEGX1_53
timestamp 1554483974
transform -1 0 1240 0 1 170
box -8 -3 104 105
use FILL  FILL_1221
timestamp 1554483974
transform 1 0 1240 0 1 170
box -8 -3 16 105
use FILL  FILL_1222
timestamp 1554483974
transform 1 0 1248 0 1 170
box -8 -3 16 105
use FILL  FILL_1223
timestamp 1554483974
transform 1 0 1256 0 1 170
box -8 -3 16 105
use FILL  FILL_1224
timestamp 1554483974
transform 1 0 1264 0 1 170
box -8 -3 16 105
use FILL  FILL_1225
timestamp 1554483974
transform 1 0 1272 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_44
timestamp 1554483974
transform 1 0 1280 0 1 170
box -8 -3 34 105
use FILL  FILL_1226
timestamp 1554483974
transform 1 0 1312 0 1 170
box -8 -3 16 105
use FILL  FILL_1227
timestamp 1554483974
transform 1 0 1320 0 1 170
box -8 -3 16 105
use FILL  FILL_1235
timestamp 1554483974
transform 1 0 1328 0 1 170
box -8 -3 16 105
use FILL  FILL_1237
timestamp 1554483974
transform 1 0 1336 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_24
timestamp 1554483974
transform -1 0 1376 0 1 170
box -8 -3 40 105
use FILL  FILL_1238
timestamp 1554483974
transform 1 0 1376 0 1 170
box -8 -3 16 105
use FILL  FILL_1239
timestamp 1554483974
transform 1 0 1384 0 1 170
box -8 -3 16 105
use FILL  FILL_1240
timestamp 1554483974
transform 1 0 1392 0 1 170
box -8 -3 16 105
use FILL  FILL_1246
timestamp 1554483974
transform 1 0 1400 0 1 170
box -8 -3 16 105
use FILL  FILL_1248
timestamp 1554483974
transform 1 0 1408 0 1 170
box -8 -3 16 105
use FILL  FILL_1250
timestamp 1554483974
transform 1 0 1416 0 1 170
box -8 -3 16 105
use FILL  FILL_1252
timestamp 1554483974
transform 1 0 1424 0 1 170
box -8 -3 16 105
use FILL  FILL_1254
timestamp 1554483974
transform 1 0 1432 0 1 170
box -8 -3 16 105
use NAND3X1  NAND3X1_25
timestamp 1554483974
transform 1 0 1440 0 1 170
box -8 -3 40 105
use FILL  FILL_1255
timestamp 1554483974
transform 1 0 1472 0 1 170
box -8 -3 16 105
use FILL  FILL_1258
timestamp 1554483974
transform 1 0 1480 0 1 170
box -8 -3 16 105
use FILL  FILL_1260
timestamp 1554483974
transform 1 0 1488 0 1 170
box -8 -3 16 105
use OAI21X1  OAI21X1_45
timestamp 1554483974
transform 1 0 1496 0 1 170
box -8 -3 34 105
use FILL  FILL_1262
timestamp 1554483974
transform 1 0 1528 0 1 170
box -8 -3 16 105
use FILL  FILL_1263
timestamp 1554483974
transform 1 0 1536 0 1 170
box -8 -3 16 105
use FILL  FILL_1264
timestamp 1554483974
transform 1 0 1544 0 1 170
box -8 -3 16 105
use FILL  FILL_1265
timestamp 1554483974
transform 1 0 1552 0 1 170
box -8 -3 16 105
use FILL  FILL_1266
timestamp 1554483974
transform 1 0 1560 0 1 170
box -8 -3 16 105
use INVX2  INVX2_84
timestamp 1554483974
transform -1 0 1584 0 1 170
box -9 -3 26 105
use FILL  FILL_1267
timestamp 1554483974
transform 1 0 1584 0 1 170
box -8 -3 16 105
use FILL  FILL_1268
timestamp 1554483974
transform 1 0 1592 0 1 170
box -8 -3 16 105
use FILL  FILL_1269
timestamp 1554483974
transform 1 0 1600 0 1 170
box -8 -3 16 105
use FILL  FILL_1270
timestamp 1554483974
transform 1 0 1608 0 1 170
box -8 -3 16 105
use NAND2X1  NAND2X1_58
timestamp 1554483974
transform 1 0 1616 0 1 170
box -8 -3 32 105
use OAI22X1  OAI22X1_25
timestamp 1554483974
transform 1 0 1640 0 1 170
box -8 -3 46 105
use DFFNEGX1  DFFNEGX1_55
timestamp 1554483974
transform 1 0 1680 0 1 170
box -8 -3 104 105
use UART_VIA1  UART_VIA1_29
timestamp 1554483974
transform 1 0 1801 0 1 170
box -10 -3 10 3
use UART_VIA1  UART_VIA1_30
timestamp 1554483974
transform 1 0 24 0 1 70
box -10 -3 10 3
use FILL  FILL_1064
timestamp 1554483974
transform 1 0 72 0 -1 170
box -8 -3 16 105
use FILL  FILL_1066
timestamp 1554483974
transform 1 0 80 0 -1 170
box -8 -3 16 105
use FILL  FILL_1068
timestamp 1554483974
transform 1 0 88 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_862
timestamp 1554483974
transform 1 0 108 0 1 115
box -3 -3 3 3
use FILL  FILL_1071
timestamp 1554483974
transform 1 0 96 0 -1 170
box -8 -3 16 105
use FILL  FILL_1072
timestamp 1554483974
transform 1 0 104 0 -1 170
box -8 -3 16 105
use FILL  FILL_1073
timestamp 1554483974
transform 1 0 112 0 -1 170
box -8 -3 16 105
use FILL  FILL_1074
timestamp 1554483974
transform 1 0 120 0 -1 170
box -8 -3 16 105
use FILL  FILL_1075
timestamp 1554483974
transform 1 0 128 0 -1 170
box -8 -3 16 105
use FILL  FILL_1076
timestamp 1554483974
transform 1 0 136 0 -1 170
box -8 -3 16 105
use FILL  FILL_1078
timestamp 1554483974
transform 1 0 144 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1166
timestamp 1554483974
transform 1 0 164 0 1 125
box -2 -2 2 2
use FILL  FILL_1083
timestamp 1554483974
transform 1 0 152 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1138
timestamp 1554483974
transform 1 0 180 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1199
timestamp 1554483974
transform 1 0 180 0 1 105
box -2 -2 2 2
use INVX2  INVX2_74
timestamp 1554483974
transform -1 0 176 0 -1 170
box -9 -3 26 105
use FILL  FILL_1084
timestamp 1554483974
transform 1 0 176 0 -1 170
box -8 -3 16 105
use FILL  FILL_1086
timestamp 1554483974
transform 1 0 184 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1167
timestamp 1554483974
transform 1 0 220 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1191
timestamp 1554483974
transform 1 0 212 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1201
timestamp 1554483974
transform 1 0 204 0 1 95
box -2 -2 2 2
use FILL  FILL_1088
timestamp 1554483974
transform 1 0 192 0 -1 170
box -8 -3 16 105
use FILL  FILL_1093
timestamp 1554483974
transform 1 0 200 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_863
timestamp 1554483974
transform 1 0 220 0 1 115
box -3 -3 3 3
use NAND3X1  NAND3X1_19
timestamp 1554483974
transform 1 0 208 0 -1 170
box -8 -3 40 105
use FILL  FILL_1094
timestamp 1554483974
transform 1 0 240 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1139
timestamp 1554483974
transform 1 0 260 0 1 135
box -2 -2 2 2
use FILL  FILL_1096
timestamp 1554483974
transform 1 0 248 0 -1 170
box -8 -3 16 105
use FILL  FILL_1097
timestamp 1554483974
transform 1 0 256 0 -1 170
box -8 -3 16 105
use FILL  FILL_1098
timestamp 1554483974
transform 1 0 264 0 -1 170
box -8 -3 16 105
use FILL  FILL_1099
timestamp 1554483974
transform 1 0 272 0 -1 170
box -8 -3 16 105
use FILL  FILL_1100
timestamp 1554483974
transform 1 0 280 0 -1 170
box -8 -3 16 105
use FILL  FILL_1101
timestamp 1554483974
transform 1 0 288 0 -1 170
box -8 -3 16 105
use FILL  FILL_1102
timestamp 1554483974
transform 1 0 296 0 -1 170
box -8 -3 16 105
use FILL  FILL_1103
timestamp 1554483974
transform 1 0 304 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1168
timestamp 1554483974
transform 1 0 332 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1192
timestamp 1554483974
transform 1 0 324 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_864
timestamp 1554483974
transform 1 0 332 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_871
timestamp 1554483974
transform 1 0 324 0 1 105
box -3 -3 3 3
use FILL  FILL_1104
timestamp 1554483974
transform 1 0 312 0 -1 170
box -8 -3 16 105
use FILL  FILL_1105
timestamp 1554483974
transform 1 0 320 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1193
timestamp 1554483974
transform 1 0 356 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_872
timestamp 1554483974
transform 1 0 356 0 1 105
box -3 -3 3 3
use OAI21X1  OAI21X1_41
timestamp 1554483974
transform 1 0 328 0 -1 170
box -8 -3 34 105
use FILL  FILL_1106
timestamp 1554483974
transform 1 0 360 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1140
timestamp 1554483974
transform 1 0 380 0 1 135
box -2 -2 2 2
use FILL  FILL_1107
timestamp 1554483974
transform 1 0 368 0 -1 170
box -8 -3 16 105
use FILL  FILL_1108
timestamp 1554483974
transform 1 0 376 0 -1 170
box -8 -3 16 105
use FILL  FILL_1109
timestamp 1554483974
transform 1 0 384 0 -1 170
box -8 -3 16 105
use FILL  FILL_1111
timestamp 1554483974
transform 1 0 392 0 -1 170
box -8 -3 16 105
use FILL  FILL_1113
timestamp 1554483974
transform 1 0 400 0 -1 170
box -8 -3 16 105
use FILL  FILL_1115
timestamp 1554483974
transform 1 0 408 0 -1 170
box -8 -3 16 105
use FILL  FILL_1117
timestamp 1554483974
transform 1 0 416 0 -1 170
box -8 -3 16 105
use FILL  FILL_1119
timestamp 1554483974
transform 1 0 424 0 -1 170
box -8 -3 16 105
use FILL  FILL_1121
timestamp 1554483974
transform 1 0 432 0 -1 170
box -8 -3 16 105
use FILL  FILL_1122
timestamp 1554483974
transform 1 0 440 0 -1 170
box -8 -3 16 105
use FILL  FILL_1123
timestamp 1554483974
transform 1 0 448 0 -1 170
box -8 -3 16 105
use FILL  FILL_1124
timestamp 1554483974
transform 1 0 456 0 -1 170
box -8 -3 16 105
use FILL  FILL_1126
timestamp 1554483974
transform 1 0 464 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1141
timestamp 1554483974
transform 1 0 484 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_850
timestamp 1554483974
transform 1 0 484 0 1 125
box -3 -3 3 3
use FILL  FILL_1128
timestamp 1554483974
transform 1 0 472 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_77
timestamp 1554483974
transform 1 0 480 0 -1 170
box -9 -3 26 105
use FILL  FILL_1132
timestamp 1554483974
transform 1 0 496 0 -1 170
box -8 -3 16 105
use FILL  FILL_1134
timestamp 1554483974
transform 1 0 504 0 -1 170
box -8 -3 16 105
use FILL  FILL_1136
timestamp 1554483974
transform 1 0 512 0 -1 170
box -8 -3 16 105
use FILL  FILL_1142
timestamp 1554483974
transform 1 0 520 0 -1 170
box -8 -3 16 105
use FILL  FILL_1143
timestamp 1554483974
transform 1 0 528 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1169
timestamp 1554483974
transform 1 0 548 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1142
timestamp 1554483974
transform 1 0 556 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_865
timestamp 1554483974
transform 1 0 548 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_851
timestamp 1554483974
transform 1 0 564 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1170
timestamp 1554483974
transform 1 0 572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1194
timestamp 1554483974
transform 1 0 556 0 1 115
box -2 -2 2 2
use FILL  FILL_1144
timestamp 1554483974
transform 1 0 536 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_866
timestamp 1554483974
transform 1 0 572 0 1 115
box -3 -3 3 3
use M3_M2  M3_M2_877
timestamp 1554483974
transform 1 0 556 0 1 95
box -3 -3 3 3
use FILL  FILL_1145
timestamp 1554483974
transform 1 0 544 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1143
timestamp 1554483974
transform 1 0 588 0 1 135
box -2 -2 2 2
use OAI21X1  OAI21X1_42
timestamp 1554483974
transform -1 0 584 0 -1 170
box -8 -3 34 105
use FILL  FILL_1146
timestamp 1554483974
transform 1 0 584 0 -1 170
box -8 -3 16 105
use FILL  FILL_1148
timestamp 1554483974
transform 1 0 592 0 -1 170
box -8 -3 16 105
use FILL  FILL_1150
timestamp 1554483974
transform 1 0 600 0 -1 170
box -8 -3 16 105
use FILL  FILL_1152
timestamp 1554483974
transform 1 0 608 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1144
timestamp 1554483974
transform 1 0 660 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_852
timestamp 1554483974
transform 1 0 636 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1171
timestamp 1554483974
transform 1 0 644 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_853
timestamp 1554483974
transform 1 0 652 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1145
timestamp 1554483974
transform 1 0 684 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1172
timestamp 1554483974
transform 1 0 676 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1195
timestamp 1554483974
transform 1 0 628 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1196
timestamp 1554483974
transform 1 0 652 0 1 115
box -2 -2 2 2
use M2_M1  M2_M1_1197
timestamp 1554483974
transform 1 0 660 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_873
timestamp 1554483974
transform 1 0 628 0 1 105
box -3 -3 3 3
use M2_M1  M2_M1_1200
timestamp 1554483974
transform 1 0 636 0 1 105
box -2 -2 2 2
use FILL  FILL_1160
timestamp 1554483974
transform 1 0 616 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_874
timestamp 1554483974
transform 1 0 660 0 1 105
box -3 -3 3 3
use M3_M2  M3_M2_878
timestamp 1554483974
transform 1 0 644 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_882
timestamp 1554483974
transform 1 0 644 0 1 85
box -3 -3 3 3
use NAND3X1  NAND3X1_21
timestamp 1554483974
transform -1 0 656 0 -1 170
box -8 -3 40 105
use M3_M2  M3_M2_854
timestamp 1554483974
transform 1 0 684 0 1 125
box -3 -3 3 3
use M3_M2  M3_M2_879
timestamp 1554483974
transform 1 0 676 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_883
timestamp 1554483974
transform 1 0 668 0 1 85
box -3 -3 3 3
use OAI21X1  OAI21X1_43
timestamp 1554483974
transform -1 0 688 0 -1 170
box -8 -3 34 105
use M2_M1  M2_M1_1146
timestamp 1554483974
transform 1 0 700 0 1 135
box -2 -2 2 2
use FILL  FILL_1161
timestamp 1554483974
transform 1 0 688 0 -1 170
box -8 -3 16 105
use FILL  FILL_1162
timestamp 1554483974
transform 1 0 696 0 -1 170
box -8 -3 16 105
use FILL  FILL_1163
timestamp 1554483974
transform 1 0 704 0 -1 170
box -8 -3 16 105
use FILL  FILL_1164
timestamp 1554483974
transform 1 0 712 0 -1 170
box -8 -3 16 105
use FILL  FILL_1165
timestamp 1554483974
transform 1 0 720 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_833
timestamp 1554483974
transform 1 0 748 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1147
timestamp 1554483974
transform 1 0 740 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1148
timestamp 1554483974
transform 1 0 748 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_855
timestamp 1554483974
transform 1 0 740 0 1 125
box -3 -3 3 3
use FILL  FILL_1167
timestamp 1554483974
transform 1 0 728 0 -1 170
box -8 -3 16 105
use FILL  FILL_1169
timestamp 1554483974
transform 1 0 736 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_834
timestamp 1554483974
transform 1 0 772 0 1 145
box -3 -3 3 3
use INVX2  INVX2_78
timestamp 1554483974
transform 1 0 744 0 -1 170
box -9 -3 26 105
use FILL  FILL_1173
timestamp 1554483974
transform 1 0 760 0 -1 170
box -8 -3 16 105
use FILL  FILL_1175
timestamp 1554483974
transform 1 0 768 0 -1 170
box -8 -3 16 105
use FILL  FILL_1177
timestamp 1554483974
transform 1 0 776 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1173
timestamp 1554483974
transform 1 0 796 0 1 125
box -2 -2 2 2
use FILL  FILL_1179
timestamp 1554483974
transform 1 0 784 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1149
timestamp 1554483974
transform 1 0 804 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_856
timestamp 1554483974
transform 1 0 804 0 1 125
box -3 -3 3 3
use FILL  FILL_1181
timestamp 1554483974
transform 1 0 792 0 -1 170
box -8 -3 16 105
use FILL  FILL_1183
timestamp 1554483974
transform 1 0 800 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1174
timestamp 1554483974
transform 1 0 820 0 1 125
box -2 -2 2 2
use INVX2  INVX2_79
timestamp 1554483974
transform 1 0 808 0 -1 170
box -9 -3 26 105
use FILL  FILL_1184
timestamp 1554483974
transform 1 0 824 0 -1 170
box -8 -3 16 105
use FILL  FILL_1185
timestamp 1554483974
transform 1 0 832 0 -1 170
box -8 -3 16 105
use FILL  FILL_1187
timestamp 1554483974
transform 1 0 840 0 -1 170
box -8 -3 16 105
use FILL  FILL_1189
timestamp 1554483974
transform 1 0 848 0 -1 170
box -8 -3 16 105
use FILL  FILL_1191
timestamp 1554483974
transform 1 0 856 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_835
timestamp 1554483974
transform 1 0 956 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1150
timestamp 1554483974
transform 1 0 956 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1175
timestamp 1554483974
transform 1 0 876 0 1 125
box -2 -2 2 2
use FILL  FILL_1201
timestamp 1554483974
transform 1 0 864 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_857
timestamp 1554483974
transform 1 0 884 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1176
timestamp 1554483974
transform 1 0 932 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_880
timestamp 1554483974
transform 1 0 892 0 1 95
box -3 -3 3 3
use M3_M2  M3_M2_881
timestamp 1554483974
transform 1 0 940 0 1 95
box -3 -3 3 3
use M2_M1  M2_M1_1151
timestamp 1554483974
transform 1 0 972 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_867
timestamp 1554483974
transform 1 0 972 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_51
timestamp 1554483974
transform -1 0 968 0 -1 170
box -8 -3 104 105
use FILL  FILL_1202
timestamp 1554483974
transform 1 0 968 0 -1 170
box -8 -3 16 105
use INVX2  INVX2_80
timestamp 1554483974
transform 1 0 976 0 -1 170
box -9 -3 26 105
use FILL  FILL_1206
timestamp 1554483974
transform 1 0 992 0 -1 170
box -8 -3 16 105
use FILL  FILL_1214
timestamp 1554483974
transform 1 0 1000 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_829
timestamp 1554483974
transform 1 0 1028 0 1 155
box -3 -3 3 3
use M3_M2  M3_M2_830
timestamp 1554483974
transform 1 0 1060 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1177
timestamp 1554483974
transform 1 0 1020 0 1 125
box -2 -2 2 2
use FILL  FILL_1215
timestamp 1554483974
transform 1 0 1008 0 -1 170
box -8 -3 16 105
use FILL  FILL_1216
timestamp 1554483974
transform 1 0 1016 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_836
timestamp 1554483974
transform 1 0 1036 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1152
timestamp 1554483974
transform 1 0 1036 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1153
timestamp 1554483974
transform 1 0 1124 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1178
timestamp 1554483974
transform 1 0 1060 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1179
timestamp 1554483974
transform 1 0 1116 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_868
timestamp 1554483974
transform 1 0 1116 0 1 115
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_52
timestamp 1554483974
transform 1 0 1024 0 -1 170
box -8 -3 104 105
use FILL  FILL_1217
timestamp 1554483974
transform 1 0 1120 0 -1 170
box -8 -3 16 105
use FILL  FILL_1219
timestamp 1554483974
transform 1 0 1128 0 -1 170
box -8 -3 16 105
use FILL  FILL_1228
timestamp 1554483974
transform 1 0 1136 0 -1 170
box -8 -3 16 105
use NOR2X1  NOR2X1_16
timestamp 1554483974
transform -1 0 1168 0 -1 170
box -8 -3 32 105
use FILL  FILL_1229
timestamp 1554483974
transform 1 0 1168 0 -1 170
box -8 -3 16 105
use FILL  FILL_1230
timestamp 1554483974
transform 1 0 1176 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1154
timestamp 1554483974
transform 1 0 1196 0 1 135
box -2 -2 2 2
use FILL  FILL_1231
timestamp 1554483974
transform 1 0 1184 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1180
timestamp 1554483974
transform 1 0 1204 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1181
timestamp 1554483974
transform 1 0 1212 0 1 125
box -2 -2 2 2
use INVX2  INVX2_81
timestamp 1554483974
transform 1 0 1192 0 -1 170
box -9 -3 26 105
use FILL  FILL_1232
timestamp 1554483974
transform 1 0 1208 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_837
timestamp 1554483974
transform 1 0 1228 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_838
timestamp 1554483974
transform 1 0 1284 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_839
timestamp 1554483974
transform 1 0 1308 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1155
timestamp 1554483974
transform 1 0 1308 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_858
timestamp 1554483974
transform 1 0 1228 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1182
timestamp 1554483974
transform 1 0 1284 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_859
timestamp 1554483974
transform 1 0 1308 0 1 125
box -3 -3 3 3
use FILL  FILL_1233
timestamp 1554483974
transform 1 0 1216 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_875
timestamp 1554483974
transform 1 0 1308 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_54
timestamp 1554483974
transform -1 0 1320 0 -1 170
box -8 -3 104 105
use FILL  FILL_1234
timestamp 1554483974
transform 1 0 1320 0 -1 170
box -8 -3 16 105
use FILL  FILL_1236
timestamp 1554483974
transform 1 0 1328 0 -1 170
box -8 -3 16 105
use FILL  FILL_1241
timestamp 1554483974
transform 1 0 1336 0 -1 170
box -8 -3 16 105
use FILL  FILL_1242
timestamp 1554483974
transform 1 0 1344 0 -1 170
box -8 -3 16 105
use FILL  FILL_1243
timestamp 1554483974
transform 1 0 1352 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_831
timestamp 1554483974
transform 1 0 1372 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1137
timestamp 1554483974
transform 1 0 1372 0 1 145
box -2 -2 2 2
use FILL  FILL_1244
timestamp 1554483974
transform 1 0 1360 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_832
timestamp 1554483974
transform 1 0 1388 0 1 155
box -3 -3 3 3
use M2_M1  M2_M1_1156
timestamp 1554483974
transform 1 0 1380 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1157
timestamp 1554483974
transform 1 0 1388 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1183
timestamp 1554483974
transform 1 0 1396 0 1 125
box -2 -2 2 2
use NOR2X1  NOR2X1_17
timestamp 1554483974
transform 1 0 1368 0 -1 170
box -8 -3 32 105
use FILL  FILL_1245
timestamp 1554483974
transform 1 0 1392 0 -1 170
box -8 -3 16 105
use FILL  FILL_1247
timestamp 1554483974
transform 1 0 1400 0 -1 170
box -8 -3 16 105
use FILL  FILL_1249
timestamp 1554483974
transform 1 0 1408 0 -1 170
box -8 -3 16 105
use FILL  FILL_1251
timestamp 1554483974
transform 1 0 1416 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1158
timestamp 1554483974
transform 1 0 1436 0 1 135
box -2 -2 2 2
use FILL  FILL_1253
timestamp 1554483974
transform 1 0 1424 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_840
timestamp 1554483974
transform 1 0 1452 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_846
timestamp 1554483974
transform 1 0 1444 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1159
timestamp 1554483974
transform 1 0 1452 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1184
timestamp 1554483974
transform 1 0 1444 0 1 125
box -2 -2 2 2
use M3_M2  M3_M2_869
timestamp 1554483974
transform 1 0 1452 0 1 115
box -3 -3 3 3
use INVX2  INVX2_82
timestamp 1554483974
transform 1 0 1432 0 -1 170
box -9 -3 26 105
use M3_M2  M3_M2_847
timestamp 1554483974
transform 1 0 1468 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1185
timestamp 1554483974
transform 1 0 1460 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1186
timestamp 1554483974
transform 1 0 1468 0 1 125
box -2 -2 2 2
use INVX2  INVX2_83
timestamp 1554483974
transform 1 0 1448 0 -1 170
box -9 -3 26 105
use FILL  FILL_1256
timestamp 1554483974
transform 1 0 1464 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_841
timestamp 1554483974
transform 1 0 1484 0 1 145
box -3 -3 3 3
use FILL  FILL_1257
timestamp 1554483974
transform 1 0 1472 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_860
timestamp 1554483974
transform 1 0 1492 0 1 125
box -3 -3 3 3
use FILL  FILL_1259
timestamp 1554483974
transform 1 0 1480 0 -1 170
box -8 -3 16 105
use FILL  FILL_1261
timestamp 1554483974
transform 1 0 1488 0 -1 170
box -8 -3 16 105
use M2_M1  M2_M1_1160
timestamp 1554483974
transform 1 0 1508 0 1 135
box -2 -2 2 2
use FILL  FILL_1271
timestamp 1554483974
transform 1 0 1496 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_842
timestamp 1554483974
transform 1 0 1532 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_843
timestamp 1554483974
transform 1 0 1572 0 1 145
box -3 -3 3 3
use M3_M2  M3_M2_844
timestamp 1554483974
transform 1 0 1620 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1161
timestamp 1554483974
transform 1 0 1532 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1162
timestamp 1554483974
transform 1 0 1620 0 1 135
box -2 -2 2 2
use M2_M1  M2_M1_1163
timestamp 1554483974
transform 1 0 1636 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_861
timestamp 1554483974
transform 1 0 1532 0 1 125
box -3 -3 3 3
use M2_M1  M2_M1_1187
timestamp 1554483974
transform 1 0 1540 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1188
timestamp 1554483974
transform 1 0 1572 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1198
timestamp 1554483974
transform 1 0 1532 0 1 115
box -2 -2 2 2
use M3_M2  M3_M2_870
timestamp 1554483974
transform 1 0 1540 0 1 115
box -3 -3 3 3
use OAI21X1  OAI21X1_46
timestamp 1554483974
transform 1 0 1504 0 -1 170
box -8 -3 34 105
use M3_M2  M3_M2_876
timestamp 1554483974
transform 1 0 1620 0 1 105
box -3 -3 3 3
use DFFNEGX1  DFFNEGX1_56
timestamp 1554483974
transform -1 0 1632 0 -1 170
box -8 -3 104 105
use M3_M2  M3_M2_848
timestamp 1554483974
transform 1 0 1660 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1164
timestamp 1554483974
transform 1 0 1668 0 1 135
box -2 -2 2 2
use INVX2  INVX2_85
timestamp 1554483974
transform 1 0 1632 0 -1 170
box -9 -3 26 105
use FILL  FILL_1272
timestamp 1554483974
transform 1 0 1648 0 -1 170
box -8 -3 16 105
use FILL  FILL_1273
timestamp 1554483974
transform 1 0 1656 0 -1 170
box -8 -3 16 105
use FILL  FILL_1274
timestamp 1554483974
transform 1 0 1664 0 -1 170
box -8 -3 16 105
use FILL  FILL_1275
timestamp 1554483974
transform 1 0 1672 0 -1 170
box -8 -3 16 105
use M3_M2  M3_M2_845
timestamp 1554483974
transform 1 0 1692 0 1 145
box -3 -3 3 3
use M2_M1  M2_M1_1165
timestamp 1554483974
transform 1 0 1692 0 1 135
box -2 -2 2 2
use M3_M2  M3_M2_849
timestamp 1554483974
transform 1 0 1716 0 1 135
box -3 -3 3 3
use M2_M1  M2_M1_1189
timestamp 1554483974
transform 1 0 1716 0 1 125
box -2 -2 2 2
use M2_M1  M2_M1_1190
timestamp 1554483974
transform 1 0 1772 0 1 125
box -2 -2 2 2
use DFFNEGX1  DFFNEGX1_57
timestamp 1554483974
transform 1 0 1680 0 -1 170
box -8 -3 104 105
use UART_VIA1  UART_VIA1_31
timestamp 1554483974
transform 1 0 1825 0 1 70
box -10 -3 10 3
use UART_VIA0  UART_VIA0_4
timestamp 1554483974
transform 1 0 48 0 1 47
box -10 -10 10 10
use UART_VIA0  UART_VIA0_5
timestamp 1554483974
transform 1 0 1801 0 1 47
box -10 -10 10 10
use UART_VIA0  UART_VIA0_6
timestamp 1554483974
transform 1 0 24 0 1 23
box -10 -10 10 10
use M3_M2  M3_M2_884
timestamp 1554483974
transform 1 0 876 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_885
timestamp 1554483974
transform 1 0 988 0 1 25
box -3 -3 3 3
use M3_M2  M3_M2_886
timestamp 1554483974
transform 1 0 420 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_887
timestamp 1554483974
transform 1 0 452 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_888
timestamp 1554483974
transform 1 0 924 0 1 15
box -3 -3 3 3
use M3_M2  M3_M2_889
timestamp 1554483974
transform 1 0 972 0 1 15
box -3 -3 3 3
use UART_VIA0  UART_VIA0_7
timestamp 1554483974
transform 1 0 1825 0 1 23
box -10 -10 10 10
<< labels >>
rlabel metal3 2 495 2 495 4 p_clka
rlabel metal3 2 825 2 825 4 p_clkb
rlabel metal2 644 1 644 1 4 p_reset
rlabel metal2 852 1638 852 1638 4 p_tx_data[7]
rlabel metal2 836 1638 836 1638 4 p_tx_data[6]
rlabel metal2 916 1638 916 1638 4 p_tx_data[5]
rlabel metal2 892 1638 892 1638 4 p_tx_data[4]
rlabel metal2 820 1638 820 1638 4 p_tx_data[3]
rlabel metal2 868 1638 868 1638 4 p_tx_data[2]
rlabel metal2 1292 1638 1292 1638 4 p_tx_data[1]
rlabel metal2 1308 1638 1308 1638 4 p_tx_data[0]
rlabel metal2 204 1 204 1 4 p_tx_rdy
rlabel metal2 564 1 564 1 4 p_rx_rdy
rlabel metal3 2 665 2 665 4 p_tx_busy
rlabel metal3 2 785 2 785 4 tx_out[7]
rlabel metal2 1020 1638 1020 1638 4 tx_out[6]
rlabel metal2 972 1638 972 1638 4 tx_out[5]
rlabel metal2 932 1638 932 1638 4 tx_out[4]
rlabel metal2 876 1 876 1 4 tx_out[3]
rlabel metal2 948 1638 948 1638 4 tx_out[2]
rlabel metal3 2 535 2 535 4 tx_out[1]
rlabel metal2 940 1 940 1 4 tx_out[0]
rlabel metal2 772 1 772 1 4 p_tx_done
rlabel metal3 2 1145 2 1145 4 tcount[3]
rlabel metal2 364 1638 364 1638 4 tcount[2]
rlabel metal2 412 1638 412 1638 4 tcount[1]
rlabel metal2 548 1638 548 1638 4 tcount[0]
rlabel metal2 452 1 452 1 4 tstate[3]
rlabel metal3 2 375 2 375 4 tstate[2]
rlabel metal3 2 415 2 415 4 tstate[1]
rlabel metal2 260 1 260 1 4 tstate[0]
rlabel metal3 2 735 2 735 4 p_tx_error
rlabel metal3 2 935 2 935 4 p_tx_idle
rlabel metal2 1196 1 1196 1 4 p_rx_busy
rlabel metal2 1356 1638 1356 1638 4 rx_out[7]
rlabel metal2 1476 1638 1476 1638 4 rx_out[6]
rlabel metal2 1452 1638 1452 1638 4 rx_out[5]
rlabel metal2 1564 1638 1564 1638 4 rx_out[4]
rlabel metal2 1548 1638 1548 1638 4 rx_out[3]
rlabel metal3 1847 1205 1847 1205 4 rx_out[2]
rlabel metal2 1228 1638 1228 1638 4 rx_out[1]
rlabel metal2 1164 1638 1164 1638 4 rx_out[0]
rlabel metal3 1847 955 1847 955 4 p_rx_done
rlabel metal2 1452 1 1452 1 4 rcount[3]
rlabel metal3 1847 475 1847 475 4 rcount[2]
rlabel metal3 1847 435 1847 435 4 rcount[1]
rlabel metal3 1847 385 1847 385 4 rcount[0]
rlabel metal2 788 1 788 1 4 rstate[3]
rlabel metal2 924 1 924 1 4 rstate[2]
rlabel metal2 756 1 756 1 4 rstate[1]
rlabel metal2 740 1 740 1 4 rstate[0]
rlabel metal3 1847 675 1847 675 4 p_rx_error
rlabel metal2 1156 1 1156 1 4 p_rx_idle
rlabel metal2 1092 1638 1092 1638 4 match
rlabel metal2 1140 1638 1140 1638 4 p_rxrxout[7]
rlabel metal2 1124 1638 1124 1638 4 p_rxrxout[6]
rlabel metal2 1204 1638 1204 1638 4 p_rxrxout[5]
rlabel metal2 1180 1638 1180 1638 4 p_rxrxout[4]
rlabel metal2 1244 1638 1244 1638 4 p_rxrxout[3]
rlabel metal2 1260 1638 1260 1638 4 p_rxrxout[2]
rlabel metal2 1276 1638 1276 1638 4 p_rxrxout[1]
rlabel metal2 1108 1638 1108 1638 4 p_rxrxout[0]
rlabel metal1 38 167 38 167 4 gnd
rlabel metal1 14 67 14 67 4 vdd
rlabel metal2 819 1632 819 1632 1 p_tx_data[3]
rlabel metal2 836 1632 836 1632 1 p_tx_data[6]
rlabel metal2 851 1632 851 1632 1 p_tx_data[7]
rlabel metal2 868 1633 868 1633 1 p_tx_data[2]
rlabel metal2 892 1633 892 1633 1 p_tx_data[4]
rlabel metal2 916 1633 916 1633 1 p_tx_data[5]
rlabel metal2 1108 1633 1108 1633 1 p_rxrxout[0]
rlabel metal2 1124 1633 1124 1633 1 p_rxrxout[6]
rlabel metal2 1140 1633 1140 1633 1 p_rxrxout[7]
rlabel metal2 1163 1633 1163 1633 1 p_rxrxout[0]
rlabel metal2 1180 1634 1180 1634 1 p_rxrxout[4]
rlabel metal2 1204 1633 1204 1633 1 p_rxrxout[5]
rlabel metal2 1243 1634 1243 1634 1 p_rxrxout[3]
rlabel metal2 1260 1635 1260 1635 5 p_rxrxout[2]
rlabel metal2 1276 1634 1276 1634 1 p_rxrxout[1]
rlabel metal2 1291 1635 1291 1635 5 p_tx_data[1]
rlabel metal2 1308 1634 1308 1634 1 p_tx_data[0]
rlabel metal3 1841 955 1841 955 1 p_rx_done
rlabel metal3 1841 674 1841 674 1 p_rx_error
rlabel metal2 1195 7 1195 7 1 p_rx_busy
rlabel metal2 1156 7 1156 7 1 p_rx_idle
rlabel metal2 772 8 772 8 1 p_tx_done
rlabel metal2 643 7 643 7 1 p_reset
rlabel metal2 564 7 564 7 1 p_rx_rdy
rlabel metal2 204 5 204 5 1 p_tx_rdy
rlabel metal3 10 664 10 664 1 p_tx_busy
rlabel metal3 10 734 10 734 1 p_tx_error
rlabel metal3 8 823 8 823 1 p_clkb
rlabel metal3 10 934 10 934 1 p_tx_idle
<< end >>
